magic
tech sky130l
timestamp 1668240734
<< m1 >>
rect 8 20 12 24
rect 8 4 12 8
<< labels >>
rlabel m1 s 8 20 12 24 6 Vdd
port 1 nsew power input
rlabel m1 s 8 4 12 8 6 GND
port 2 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 16 28
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
