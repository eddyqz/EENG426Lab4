magic
tech sky130l
timestamp 1668327008
<< ndiffusion >>
rect 8 13 13 16
rect 8 10 9 13
rect 12 10 13 13
rect 8 6 13 10
rect 15 6 20 16
rect 22 13 27 16
rect 22 10 23 13
rect 26 10 27 13
rect 22 6 27 10
<< ndc >>
rect 9 10 12 13
rect 23 10 26 13
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 30 13 31
rect 8 27 9 30
rect 12 27 13 30
rect 8 23 13 27
rect 15 27 20 31
rect 15 24 16 27
rect 19 24 20 27
rect 15 23 20 24
rect 22 30 27 31
rect 22 27 23 30
rect 26 27 27 30
rect 22 23 27 27
<< pdc >>
rect 9 27 12 30
rect 16 24 19 27
rect 23 27 26 30
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
<< polysilicon >>
rect 13 31 15 33
rect 20 31 22 33
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 10 3 15 4
rect 10 0 11 3
rect 14 0 15 3
rect 10 -1 15 0
rect 20 4 22 6
rect 20 3 25 4
rect 20 0 21 3
rect 24 0 25 3
rect 20 -1 25 0
<< pc >>
rect 11 0 14 3
rect 21 0 24 3
<< m1 >>
rect 8 36 13 41
rect 22 36 27 41
rect 9 31 12 36
rect 23 31 26 36
rect 8 30 13 31
rect 8 27 9 30
rect 12 27 13 30
rect 22 30 27 31
rect 8 26 13 27
rect 16 27 19 28
rect 22 27 23 30
rect 26 27 27 30
rect 22 26 27 27
rect 16 21 19 24
rect 16 18 33 21
rect 3 13 13 14
rect 3 10 4 13
rect 7 10 9 13
rect 12 10 13 13
rect 3 9 13 10
rect 22 13 27 14
rect 30 13 33 18
rect 22 10 23 13
rect 26 10 33 13
rect 22 9 27 10
rect 10 3 15 4
rect 10 0 11 3
rect 14 0 15 3
rect 10 -1 15 0
rect 20 3 25 4
rect 20 0 21 3
rect 24 0 25 3
rect 20 -1 25 0
<< m2c >>
rect 4 10 7 13
<< m2 >>
rect 8 40 13 41
rect 22 40 27 41
rect 8 37 27 40
rect 8 36 13 37
rect 22 36 27 37
rect 1 13 8 14
rect 1 10 4 13
rect 7 10 8 13
rect 1 9 8 10
<< labels >>
rlabel ndiffusion 23 7 23 7 3 Y
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 B
rlabel polysilicon 21 22 21 22 3 B
rlabel pdiffusion 16 24 16 24 3 Y
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m2 14 39 14 39 5 Vdd
rlabel m1 31 19 31 19 7 Y
rlabel m2 2 11 2 11 3 GND
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 40 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
