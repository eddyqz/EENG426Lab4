magic
tech sky130l
timestamp 1668540001
<< ndiffusion >>
rect 16 26 21 28
rect 16 23 17 26
rect 20 23 21 26
rect 16 22 21 23
rect 23 26 29 28
rect 23 23 25 26
rect 28 23 29 26
rect 23 22 29 23
<< ndc >>
rect 17 23 20 26
rect 25 23 28 26
<< ntransistor >>
rect 21 22 23 28
<< pdiffusion >>
rect 14 40 20 43
rect 14 37 15 40
rect 18 37 20 40
rect 14 35 20 37
rect 24 39 29 43
rect 24 36 25 39
rect 28 36 29 39
rect 24 35 29 36
<< pdc >>
rect 15 37 18 40
rect 25 36 28 39
<< ptransistor >>
rect 20 35 24 43
<< polysilicon >>
rect 20 43 24 45
rect 5 34 10 35
rect 20 34 24 35
rect 5 31 6 34
rect 9 31 24 34
rect 5 30 24 31
rect 21 28 23 30
rect 21 20 23 22
<< pc >>
rect 6 31 9 34
<< m1 >>
rect 16 47 20 61
rect 6 44 20 47
rect 24 48 29 61
rect 24 45 25 48
rect 28 45 29 48
rect 24 44 29 45
rect 32 45 36 48
rect 32 44 39 45
rect 6 35 9 44
rect 33 41 35 44
rect 38 41 39 44
rect 14 40 19 41
rect 14 37 15 40
rect 18 37 19 40
rect 14 36 19 37
rect 25 39 28 41
rect 33 39 39 41
rect 28 36 29 39
rect 5 34 10 35
rect 5 31 6 34
rect 9 31 10 34
rect 5 30 10 31
rect 25 27 28 36
rect 16 26 21 27
rect 16 23 17 26
rect 20 23 21 26
rect 16 22 21 23
rect 24 26 30 27
rect 24 23 25 26
rect 28 23 30 26
rect 24 22 30 23
rect 16 16 20 22
rect 33 16 36 39
rect 16 13 36 16
rect 24 9 29 10
rect 24 6 25 9
rect 28 6 29 9
rect 24 5 29 6
<< m2c >>
rect 25 45 28 48
rect 35 41 38 44
rect 15 37 18 40
rect 25 23 28 26
rect 25 6 28 9
<< m2 >>
rect 16 53 28 56
rect 16 41 20 53
rect 25 49 28 53
rect 24 48 29 49
rect 24 45 25 48
rect 28 45 29 48
rect 24 44 29 45
rect 33 44 39 45
rect 14 40 20 41
rect 14 37 15 40
rect 18 37 20 40
rect 33 41 35 44
rect 38 41 39 44
rect 33 39 39 41
rect 14 36 19 37
rect 24 26 29 27
rect 24 23 25 26
rect 28 23 29 26
rect 24 9 29 23
rect 24 6 25 9
rect 28 6 29 9
rect 24 5 29 6
<< labels >>
rlabel polysilicon 22 29 22 29 3 A
rlabel polysilicon 21 35 21 35 3 A
rlabel ndiffusion 24 23 24 23 3 Y
rlabel ndiffusion 24 24 24 24 3 Y
rlabel ndiffusion 24 27 24 27 3 Y
rlabel pdiffusion 25 36 25 36 3 Y
rlabel pdiffusion 25 37 25 37 3 Y
rlabel pdiffusion 25 40 25 40 3 Y
rlabel polysilicon 21 44 21 44 3 A
rlabel polysilicon 22 21 22 21 3 A
rlabel ntransistor 22 23 22 23 3 A
rlabel ptransistor 21 36 21 36 3 A
rlabel pdiffusion 15 36 15 36 3 Vdd
rlabel m1 29 37 29 37 3 Y
port 1 e
rlabel m1 33 45 33 45 3 GND
rlabel m1 26 28 26 28 3 Y
port 1 e
rlabel pdc 26 37 26 37 3 Y
port 1 e
rlabel m1 26 40 26 40 3 Y
port 1 e
rlabel m1 25 23 25 23 3 Y
port 1 e
rlabel m1 17 48 17 48 3 A
port 2 e
rlabel m1 10 32 10 32 3 A
port 2 e
rlabel pc 7 32 7 32 3 A
port 2 e
rlabel m1 7 36 7 36 3 A
port 2 e
rlabel m1 7 45 7 45 3 A
port 2 e
rlabel m1 6 31 6 31 3 A
port 2 e
rlabel m1 6 32 6 32 3 A
port 2 e
rlabel m1 6 35 6 35 3 A
port 2 e
rlabel m2 29 46 29 46 3 Vdd
rlabel m2c 26 46 26 46 3 Vdd
rlabel m2 26 50 26 50 3 Vdd
rlabel m2 29 7 29 7 3 Y
port 1 e
rlabel m2 29 24 29 24 3 Y
port 1 e
rlabel m2 25 45 25 45 3 Vdd
rlabel m2 25 46 25 46 3 Vdd
rlabel m2 25 49 25 49 3 Vdd
rlabel m2c 26 7 26 7 3 Y
port 1 e
rlabel m2c 26 24 26 24 3 Y
port 1 e
rlabel m2 25 6 25 6 3 Y
port 1 e
rlabel m2 25 7 25 7 3 Y
port 1 e
rlabel m2 25 10 25 10 3 Y
port 1 e
rlabel m2 25 24 25 24 3 Y
port 1 e
rlabel m2 25 27 25 27 3 Y
port 1 e
rlabel m2 19 38 19 38 3 Vdd
rlabel m2 17 42 17 42 3 Vdd
rlabel m2 17 54 17 54 3 Vdd
rlabel m2c 16 38 16 38 3 Vdd
rlabel m2 15 37 15 37 3 Vdd
rlabel m2 15 38 15 38 3 Vdd
rlabel m2 15 41 15 41 3 Vdd
rlabel m2c 36 42 36 42 7 GND
rlabel ndc 18 24 18 24 1 GND
rlabel m1 18 18 18 18 1 GND
<< end >>
