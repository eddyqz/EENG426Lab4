magic
tech sky130l
timestamp 1668469005
<< checkpaint >>
rect -26 28 68 98
rect -25 26 68 28
rect -24 -19 68 26
rect -24 -22 59 -19
rect -24 -24 54 -22
rect -24 -28 51 -24
rect -24 -29 44 -28
<< ndiffusion >>
rect 8 17 13 20
rect 8 14 9 17
rect 12 14 13 17
rect 8 10 13 14
rect 15 17 20 20
rect 15 14 16 17
rect 19 14 20 17
rect 15 10 20 14
rect 22 17 27 20
rect 22 14 23 17
rect 26 14 27 17
rect 22 10 27 14
<< ndc >>
rect 9 14 12 17
rect 16 14 19 17
rect 23 14 26 17
<< ntransistor >>
rect 13 10 15 20
rect 20 10 22 20
<< pdiffusion >>
rect 8 43 13 57
rect 8 40 9 43
rect 12 40 13 43
rect 8 27 13 40
rect 15 27 20 57
rect 22 33 27 57
rect 22 30 23 33
rect 26 30 27 33
rect 22 27 27 30
<< pdc >>
rect 9 40 12 43
rect 23 30 26 33
<< ptransistor >>
rect 13 27 15 57
rect 20 27 22 57
<< polysilicon >>
rect 6 64 11 65
rect 6 61 7 64
rect 10 61 11 64
rect 6 60 11 61
rect 18 64 23 65
rect 18 61 19 64
rect 22 61 23 64
rect 18 60 23 61
rect 7 58 15 60
rect 13 57 15 58
rect 20 57 22 60
rect 13 20 15 27
rect 20 20 22 27
rect 13 8 15 10
rect 20 8 22 10
<< pc >>
rect 7 61 10 64
rect 19 61 22 64
<< m1 >>
rect 6 64 11 66
rect 6 61 7 64
rect 10 61 11 64
rect 6 60 11 61
rect 18 64 23 66
rect 18 61 19 64
rect 22 61 23 64
rect 18 60 23 61
rect 26 45 30 66
rect 8 43 13 44
rect 8 40 9 43
rect 12 40 13 43
rect 8 39 13 40
rect 25 43 30 45
rect 25 40 26 43
rect 29 40 30 43
rect 25 39 30 40
rect 23 33 26 34
rect 23 25 26 30
rect 16 22 26 25
rect 8 17 13 18
rect 8 14 9 17
rect 12 14 13 17
rect 8 13 13 14
rect 16 17 19 22
rect 33 18 36 66
rect 16 7 19 14
rect 22 17 36 18
rect 22 14 23 17
rect 26 14 36 17
rect 22 13 36 14
rect 8 4 19 7
rect 8 3 12 4
<< m2c >>
rect 9 40 12 43
rect 26 40 29 43
rect 9 14 12 17
rect 23 14 26 17
<< m2 >>
rect 8 43 30 44
rect 8 40 9 43
rect 12 40 26 43
rect 29 40 30 43
rect 8 39 30 40
rect 8 17 27 18
rect 8 14 9 17
rect 12 14 23 17
rect 26 14 27 17
rect 8 13 27 14
<< labels >>
rlabel pdiffusion 27 31 27 31 3 Y
rlabel polysilicon 21 58 21 58 3 B
rlabel ndiffusion 23 11 23 11 3 GND
rlabel ndiffusion 20 15 20 15 3 Y
rlabel pdiffusion 23 28 23 28 3 Y
rlabel pdiffusion 23 31 23 31 3 Y
rlabel pdiffusion 23 34 23 34 3 Y
rlabel polysilicon 21 9 21 9 3 B
rlabel ntransistor 21 11 21 11 3 B
rlabel polysilicon 21 21 21 21 3 B
rlabel ptransistor 21 28 21 28 3 B
rlabel ndiffusion 16 11 16 11 3 Y
rlabel ndiffusion 16 15 16 15 3 Y
rlabel ndiffusion 16 18 16 18 3 Y
rlabel polysilicon 14 58 14 58 3 A
rlabel polysilicon 14 9 14 9 3 A
rlabel ntransistor 14 11 14 11 3 A
rlabel polysilicon 14 21 14 21 3 A
rlabel ptransistor 14 28 14 28 3 A
rlabel ndiffusion 9 11 9 11 3 GND
rlabel pdiffusion 9 28 9 28 3 Vdd
rlabel polysilicon 8 59 8 59 3 A
rlabel m1 34 19 34 19 3 GND
rlabel m1 27 46 27 46 3 Vdd
rlabel m1 23 15 23 15 3 GND
rlabel m1 23 18 23 18 3 GND
rlabel m1 26 40 26 40 3 Vdd
rlabel m1 26 41 26 41 3 Vdd
rlabel m1 26 44 26 44 3 Vdd
rlabel m1 24 26 24 26 3 Y
port 1 e
rlabel pdc 24 31 24 31 3 Y
port 1 e
rlabel m1 24 34 24 34 3 Y
port 1 e
rlabel m1 23 62 23 62 3 B
port 2 e
rlabel m1 23 14 23 14 3 GND
rlabel ndc 17 15 17 15 3 Y
port 1 e
rlabel pc 20 62 20 62 3 B
port 2 e
rlabel m1 19 61 19 61 3 B
port 2 e
rlabel m1 19 62 19 62 3 B
port 2 e
rlabel m1 19 65 19 65 3 B
port 2 e
rlabel m1 17 8 17 8 3 Y
port 1 e
rlabel m1 17 18 17 18 3 Y
port 1 e
rlabel m1 17 23 17 23 3 Y
port 1 e
rlabel m1 9 4 9 4 3 Y
port 1 e
rlabel m1 9 5 9 5 3 Y
port 1 e
rlabel m1 11 62 11 62 3 A
port 3 e
rlabel pc 8 62 8 62 3 A
port 3 e
rlabel m1 7 61 7 61 3 A
port 3 e
rlabel m1 7 62 7 62 3 A
port 3 e
rlabel m1 7 65 7 65 3 A
port 3 e
rlabel m2 27 15 27 15 3 GND
rlabel m2 30 41 30 41 3 Vdd
rlabel m2c 24 15 24 15 3 GND
rlabel m2c 27 41 27 41 3 Vdd
rlabel m2 13 15 13 15 3 GND
rlabel m2 13 41 13 41 3 Vdd
rlabel m2c 10 15 10 15 3 GND
rlabel m2c 10 41 10 41 3 Vdd
rlabel m2 9 14 9 14 3 GND
rlabel m2 9 15 9 15 3 GND
rlabel m2 9 18 9 18 3 GND
rlabel m2 9 40 9 40 3 Vdd
rlabel m2 9 41 9 41 3 Vdd
rlabel m2 9 44 9 44 3 Vdd
<< end >>
