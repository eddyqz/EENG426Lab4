magic
tech sky130l
timestamp 1668327500
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 24 13 34
rect 8 21 9 24
rect 12 21 13 24
rect 8 19 13 21
rect 15 19 20 34
rect 22 24 27 34
rect 22 21 23 24
rect 26 21 27 24
rect 22 19 27 21
<< pdc >>
rect 9 21 12 24
rect 23 21 26 24
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 8 42 15 43
rect 8 39 9 42
rect 12 39 15 42
rect 8 38 15 39
rect 13 34 15 38
rect 20 42 27 43
rect 20 39 23 42
rect 26 39 27 42
rect 20 38 27 39
rect 20 34 22 38
rect 13 12 15 19
rect 20 12 22 19
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 9 39 12 42
rect 23 39 26 42
<< m1 >>
rect 8 42 13 43
rect 8 39 9 42
rect 12 39 13 42
rect 8 38 13 39
rect 22 42 27 43
rect 22 39 23 42
rect 26 39 27 42
rect 22 38 27 39
rect 3 24 13 25
rect 3 21 4 24
rect 7 21 9 24
rect 12 21 13 24
rect 3 20 13 21
rect 22 24 27 25
rect 22 21 23 24
rect 26 21 27 24
rect 22 20 27 21
rect 23 17 26 20
rect 16 14 26 17
rect 9 10 12 11
rect 9 4 12 7
rect 16 10 19 14
rect 16 6 19 7
rect 23 10 26 11
rect 23 4 26 7
rect 8 3 13 4
rect 8 0 9 3
rect 12 0 13 3
rect 8 -1 13 0
rect 22 3 27 4
rect 22 0 23 3
rect 26 0 27 3
rect 22 -1 27 0
<< m2c >>
rect 4 21 7 24
rect 9 0 12 3
rect 23 0 26 3
<< m2 >>
rect 1 24 8 25
rect 1 21 4 24
rect 7 21 8 24
rect 1 20 8 21
rect 8 3 13 4
rect 22 3 27 4
rect 8 0 9 3
rect 12 0 23 3
rect 26 0 27 3
rect 8 -1 13 0
rect 22 -1 27 0
<< labels >>
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Y
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m2 17 1 17 1 1 GND
rlabel m1 18 15 18 15 1 Y
rlabel m2 2 22 2 22 3 Vdd
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 40 44
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
