magic
tech sky130l
timestamp 1668469005
<< checkpaint >>
rect -10 145 91 148
rect -10 132 109 145
rect -18 97 115 132
rect -18 64 139 97
rect -19 49 139 64
rect -23 27 139 49
rect -23 -19 138 27
rect -19 -29 138 -19
<< ndiffusion >>
rect 23 31 29 36
rect 23 28 24 31
rect 27 28 29 31
rect 23 26 29 28
rect 31 26 36 36
rect 38 31 43 36
rect 38 28 39 31
rect 42 28 43 31
rect 49 34 55 36
rect 49 31 50 34
rect 53 31 55 34
rect 49 30 55 31
rect 57 30 64 36
rect 38 26 43 28
rect 58 27 59 30
rect 62 27 64 30
rect 58 26 64 27
rect 66 31 72 36
rect 66 28 68 31
rect 71 28 72 31
rect 66 26 72 28
rect 78 35 83 36
rect 78 32 79 35
rect 82 32 83 35
rect 78 26 83 32
rect 85 33 93 36
rect 85 30 89 33
rect 92 30 93 33
rect 85 26 93 30
<< ndc >>
rect 24 28 27 31
rect 39 28 42 31
rect 50 31 53 34
rect 59 27 62 30
rect 68 28 71 31
rect 79 32 82 35
rect 89 30 92 33
<< ntransistor >>
rect 29 26 31 36
rect 36 26 38 36
rect 55 30 57 36
rect 64 26 66 36
rect 83 26 85 36
<< pdiffusion >>
rect 21 53 29 58
rect 20 52 29 53
rect 20 48 21 52
rect 25 48 29 52
rect 20 47 29 48
rect 21 43 29 47
rect 31 51 35 58
rect 31 50 36 51
rect 31 47 32 50
rect 35 47 36 50
rect 31 43 36 47
rect 38 50 44 51
rect 38 47 40 50
rect 43 47 44 50
rect 38 43 44 47
rect 50 48 55 58
rect 50 45 51 48
rect 54 45 55 48
rect 50 43 55 45
rect 57 43 64 58
rect 66 56 71 58
rect 66 53 67 56
rect 70 53 71 56
rect 66 43 71 53
rect 78 49 83 58
rect 77 48 83 49
rect 77 45 79 48
rect 82 45 83 48
rect 77 43 83 45
rect 85 52 92 58
rect 85 49 88 52
rect 91 49 92 52
rect 85 43 92 49
<< pdc >>
rect 21 48 25 52
rect 32 47 35 50
rect 40 47 43 50
rect 51 45 54 48
rect 67 53 70 56
rect 79 45 82 48
rect 88 49 91 52
<< ptransistor >>
rect 29 43 31 58
rect 36 43 38 51
rect 55 43 57 58
rect 64 43 66 58
rect 83 43 85 58
<< polysilicon >>
rect 61 85 67 86
rect 61 81 62 85
rect 66 81 67 85
rect 61 80 67 81
rect 53 68 59 69
rect 22 66 28 67
rect 22 62 23 66
rect 27 62 28 66
rect 53 65 54 68
rect 52 64 54 65
rect 58 64 59 68
rect 52 63 59 64
rect 52 62 57 63
rect 22 61 28 62
rect 23 59 31 61
rect 29 58 31 59
rect 46 60 57 62
rect 46 55 48 60
rect 55 58 57 60
rect 64 58 66 80
rect 83 58 85 60
rect 36 53 48 55
rect 36 51 38 53
rect 29 36 31 43
rect 36 36 38 43
rect 55 36 57 43
rect 64 36 66 43
rect 83 36 85 43
rect 55 28 57 30
rect 29 24 31 26
rect 36 24 38 26
rect 64 24 66 26
rect 83 16 85 26
rect 81 15 87 16
rect 81 11 82 15
rect 86 11 87 15
rect 81 10 87 11
<< pc >>
rect 62 81 66 85
rect 23 62 27 66
rect 54 64 58 68
rect 82 11 86 15
<< m1 >>
rect 22 115 28 116
rect 22 111 23 115
rect 27 111 28 115
rect 40 115 45 116
rect 40 112 41 115
rect 44 112 45 115
rect 40 111 45 112
rect 53 115 59 116
rect 53 111 54 115
rect 58 111 59 115
rect 22 110 28 111
rect 53 110 59 111
rect 71 112 77 113
rect 71 108 72 112
rect 76 108 77 112
rect 71 107 77 108
rect 14 97 83 100
rect 14 51 17 97
rect 32 91 76 94
rect 22 66 28 67
rect 22 62 23 66
rect 27 62 28 66
rect 22 61 28 62
rect 24 60 28 61
rect 20 52 26 53
rect 20 51 21 52
rect 14 48 21 51
rect 25 48 26 52
rect 20 47 26 48
rect 32 50 35 91
rect 61 85 67 86
rect 40 81 62 85
rect 66 81 67 85
rect 72 82 76 87
rect 40 64 44 81
rect 61 80 67 81
rect 40 61 41 64
rect 53 68 59 69
rect 53 64 54 68
rect 58 64 59 68
rect 73 64 76 82
rect 80 64 83 97
rect 101 64 107 65
rect 53 63 60 64
rect 40 60 44 61
rect 56 60 60 63
rect 68 60 76 64
rect 79 61 83 64
rect 68 57 71 60
rect 66 56 71 57
rect 66 53 67 56
rect 70 53 71 56
rect 66 52 71 53
rect 32 46 35 47
rect 40 50 43 51
rect 79 49 82 61
rect 88 60 102 64
rect 106 60 107 64
rect 101 59 107 60
rect 87 52 92 53
rect 87 49 88 52
rect 91 49 92 52
rect 50 48 55 49
rect 40 46 43 47
rect 46 45 51 48
rect 54 45 55 48
rect 46 44 55 45
rect 78 48 83 49
rect 87 48 92 49
rect 78 45 79 48
rect 82 45 83 48
rect 78 44 83 45
rect 46 41 49 44
rect 44 40 49 41
rect 41 38 49 40
rect 41 37 47 38
rect 41 32 44 37
rect 78 35 83 36
rect 50 34 53 35
rect 23 31 28 32
rect 23 28 24 31
rect 27 28 28 31
rect 23 27 28 28
rect 38 31 44 32
rect 49 31 50 34
rect 78 32 79 35
rect 82 32 83 35
rect 67 31 71 32
rect 78 31 83 32
rect 88 33 93 34
rect 38 28 39 31
rect 42 29 44 31
rect 42 28 43 29
rect 38 27 43 28
rect 40 17 43 27
rect 9 14 43 17
rect 50 16 53 31
rect 58 30 63 31
rect 58 27 59 30
rect 62 27 63 30
rect 67 28 68 31
rect 71 28 72 31
rect 88 30 89 33
rect 92 30 93 33
rect 88 29 93 30
rect 67 27 72 28
rect 58 26 63 27
rect 48 15 53 16
rect 81 15 87 16
rect 9 13 25 14
rect 48 12 49 15
rect 52 12 82 15
rect 48 11 53 12
rect 81 11 82 12
rect 86 11 87 15
rect 81 10 87 11
<< m2c >>
rect 23 111 27 115
rect 41 112 44 115
rect 54 111 58 115
rect 72 108 76 112
rect 23 62 27 66
rect 72 87 76 91
rect 41 61 44 64
rect 54 64 58 68
rect 40 47 43 50
rect 102 60 106 64
rect 88 49 91 52
rect 51 45 54 48
rect 24 28 27 31
rect 79 32 82 35
rect 59 27 62 30
rect 68 28 71 31
rect 89 30 92 33
rect 49 12 52 15
<< m2 >>
rect 22 115 28 116
rect 22 111 23 115
rect 27 111 28 115
rect 22 66 28 111
rect 22 62 23 66
rect 27 62 28 66
rect 22 61 28 62
rect 40 115 45 116
rect 40 112 41 115
rect 44 112 45 115
rect 40 64 45 112
rect 40 61 41 64
rect 44 61 45 64
rect 53 115 59 116
rect 53 111 54 115
rect 58 111 59 115
rect 53 68 59 111
rect 71 112 77 113
rect 71 108 72 112
rect 76 108 77 112
rect 71 91 77 108
rect 71 87 72 91
rect 76 87 77 91
rect 71 86 77 87
rect 53 64 54 68
rect 58 64 59 68
rect 53 63 59 64
rect 101 64 107 65
rect 40 60 45 61
rect 101 60 102 64
rect 106 60 107 64
rect 101 59 107 60
rect 51 53 57 54
rect 51 52 92 53
rect 51 51 88 52
rect 39 50 44 51
rect 39 47 40 50
rect 43 47 44 50
rect 51 49 54 51
rect 57 50 88 51
rect 87 49 88 50
rect 91 49 92 52
rect 39 46 44 47
rect 13 31 28 32
rect 13 28 24 31
rect 27 28 28 31
rect 13 6 17 28
rect 23 27 28 28
rect 41 16 44 46
rect 50 48 55 49
rect 87 48 92 49
rect 50 45 51 48
rect 54 45 55 48
rect 50 44 55 45
rect 89 41 91 48
rect 79 39 91 41
rect 79 36 82 39
rect 78 35 83 36
rect 78 32 79 35
rect 82 32 83 35
rect 67 31 72 32
rect 78 31 83 32
rect 88 33 93 34
rect 88 31 89 33
rect 58 30 63 31
rect 58 27 59 30
rect 62 27 63 30
rect 67 28 68 31
rect 71 30 89 31
rect 92 30 93 33
rect 71 29 93 30
rect 71 28 72 29
rect 67 27 72 28
rect 58 26 63 27
rect 41 15 53 16
rect 41 12 49 15
rect 52 12 53 15
rect 48 11 53 12
rect 59 6 62 26
rect 102 6 106 59
rect 13 3 106 6
<< labels >>
rlabel polysilicon 65 59 65 59 3 B
rlabel polysilicon 62 82 62 82 3 B
rlabel ndiffusion 86 27 86 27 3 #10
rlabel ndiffusion 86 31 86 31 3 #10
rlabel ndiffusion 86 34 86 34 3 #10
rlabel polysilicon 84 37 84 37 3 _S
rlabel pdiffusion 86 44 86 44 3 Y
rlabel pdiffusion 86 50 86 50 3 Y
rlabel pdiffusion 86 53 86 53 3 Y
rlabel polysilicon 84 59 84 59 3 _S
rlabel ntransistor 84 27 84 27 3 _S
rlabel ptransistor 84 44 84 44 3 _S
rlabel pdiffusion 79 50 79 50 3 #5
rlabel pdiffusion 67 44 67 44 3 Vdd
rlabel polysilicon 54 66 54 66 3 S
rlabel ndiffusion 79 27 79 27 3 Y
rlabel pdiffusion 78 44 78 44 3 #5
rlabel pdiffusion 78 46 78 46 3 #5
rlabel pdiffusion 78 49 78 49 3 #5
rlabel ndiffusion 58 31 58 31 3 GND
rlabel polysilicon 65 37 65 37 3 B
rlabel ptransistor 65 44 65 44 3 B
rlabel polysilicon 56 59 56 59 3 S
rlabel polysilicon 53 63 53 63 3 S
rlabel polysilicon 53 64 53 64 3 S
rlabel polysilicon 53 65 53 65 3 S
rlabel polysilicon 56 29 56 29 3 S
rlabel ntransistor 56 31 56 31 3 S
rlabel ndiffusion 67 27 67 27 3 #10
rlabel ndiffusion 67 29 67 29 3 #10
rlabel ndiffusion 67 32 67 32 3 #10
rlabel ndiffusion 50 31 50 31 3 _S
rlabel ndiffusion 54 32 54 32 3 _S
rlabel polysilicon 56 37 56 37 3 S
rlabel ptransistor 56 44 56 44 3 S
rlabel ntransistor 65 27 65 27 3 B
rlabel pdiffusion 51 44 51 44 3 Y
rlabel polysilicon 47 56 47 56 3 S
rlabel polysilicon 47 61 47 61 3 S
rlabel ndiffusion 50 35 50 35 3 _S
rlabel polysilicon 65 25 65 25 3 B
rlabel ndiffusion 39 27 39 27 3 Y
rlabel polysilicon 37 37 37 37 3 S
rlabel polysilicon 84 17 84 17 3 _S
rlabel polysilicon 37 25 37 25 3 S
rlabel ntransistor 37 27 37 27 3 S
rlabel pdiffusion 39 44 39 44 3 _S
rlabel pdiffusion 39 48 39 48 3 _S
rlabel pdiffusion 39 51 39 51 3 _S
rlabel pdiffusion 36 48 36 48 3 Vdd
rlabel polysilicon 37 52 37 52 3 S
rlabel polysilicon 37 54 37 54 3 S
rlabel polysilicon 30 59 30 59 3 A
rlabel polysilicon 30 37 30 37 3 A
rlabel ptransistor 37 44 37 44 3 S
rlabel polysilicon 30 25 30 25 3 A
rlabel ntransistor 30 27 30 27 3 A
rlabel pdiffusion 32 44 32 44 3 Vdd
rlabel pdiffusion 32 48 32 48 3 Vdd
rlabel pdiffusion 32 51 32 51 3 Vdd
rlabel pdiffusion 32 52 32 52 3 Vdd
rlabel polysilicon 24 60 24 60 3 A
rlabel ndiffusion 24 27 24 27 3 GND
rlabel ptransistor 30 44 30 44 3 A
rlabel pdiffusion 22 44 22 44 3 #5
rlabel pdiffusion 22 54 22 54 3 #5
rlabel pdiffusion 21 49 21 49 3 #5
rlabel m1 81 65 81 65 3 #5
rlabel m1 74 65 74 65 3 Vdd
rlabel m1 89 61 89 61 3 GND
rlabel m1 73 83 73 83 3 Vdd
rlabel m1 83 46 83 46 3 #5
rlabel m1 88 53 88 53 3 Y
port 1 e
rlabel m1 80 62 80 62 3 #5
rlabel pdc 80 46 80 46 3 #5
rlabel m1 80 50 80 50 3 #5
rlabel m1 72 108 72 108 3 Vdd
rlabel m1 79 46 79 46 3 #5
rlabel m1 79 49 79 49 3 #5
rlabel m1 71 54 71 54 3 Vdd
rlabel m1 69 58 69 58 3 Vdd
rlabel m1 69 61 69 61 3 Vdd
rlabel pdc 68 54 68 54 3 Vdd
rlabel m1 67 53 67 53 3 Vdd
rlabel m1 67 54 67 54 3 Vdd
rlabel m1 67 57 67 57 3 Vdd
rlabel m1 62 86 62 86 3 B
port 2 e
rlabel m1 62 81 62 81 3 B
port 2 e
rlabel m1 79 45 79 45 3 #5
rlabel m1 57 61 57 61 3 S
port 3 e
rlabel m1 54 111 54 111 3 S
port 3 e
rlabel ndc 51 32 51 32 3 _S
rlabel m1 51 35 51 35 3 _S
rlabel m1 50 32 50 32 3 _S
rlabel m1 47 42 47 42 3 Y
port 1 e
rlabel m1 47 45 47 45 3 Y
port 1 e
rlabel m1 47 46 47 46 3 Y
port 1 e
rlabel m1 45 41 45 41 3 Y
port 1 e
rlabel m1 89 30 89 30 3 #10
rlabel m1 89 31 89 31 3 #10
rlabel m1 67 82 67 82 3 B
port 2 e
rlabel m1 42 33 42 33 3 Y
port 1 e
rlabel m1 42 38 42 38 3 Y
port 1 e
rlabel m1 42 39 42 39 3 Y
port 1 e
rlabel pc 63 82 63 82 3 B
port 2 e
rlabel m1 87 12 87 12 3 _S
rlabel m1 43 29 43 29 3 Y
port 1 e
rlabel m1 43 30 43 30 3 Y
port 1 e
rlabel m1 41 47 41 47 3 _S
rlabel m1 41 51 41 51 3 _S
rlabel m1 41 82 41 82 3 B
port 2 e
rlabel m1 41 112 41 112 3 B
port 2 e
rlabel pc 83 12 83 12 3 _S
rlabel ndc 40 29 40 29 3 Y
port 1 e
rlabel m1 82 11 82 11 3 _S
rlabel m1 82 12 82 12 3 _S
rlabel m1 39 29 39 29 3 Y
port 1 e
rlabel m1 39 32 39 32 3 Y
port 1 e
rlabel m1 49 13 49 13 3 _S
rlabel m1 25 61 25 61 3 A
port 4 e
rlabel m1 33 92 33 92 3 Vdd
rlabel m1 41 18 41 18 3 Y
port 1 e
rlabel m1 39 28 39 28 3 Y
port 1 e
rlabel m1 33 47 33 47 3 Vdd
rlabel pdc 33 48 33 48 3 Vdd
rlabel m1 33 51 33 51 3 Vdd
rlabel m1 82 16 82 16 3 _S
rlabel m1 24 29 24 29 3 GND
rlabel m1 24 32 24 32 3 GND
rlabel m1 51 17 51 17 3 _S
rlabel m1 26 49 26 49 3 #5
rlabel m1 21 52 21 52 3 #5
rlabel m1 21 53 21 53 3 #5
rlabel m1 23 111 23 111 3 A
port 4 e
rlabel m1 49 16 49 16 3 _S
rlabel m1 21 48 21 48 3 #5
rlabel pdc 22 49 22 49 3 #5
rlabel m1 15 49 15 49 3 #5
rlabel m1 15 52 15 52 3 #5
rlabel m1 15 98 15 98 3 #5
rlabel m1 10 14 10 14 3 Y
port 1 e
rlabel m1 10 15 10 15 3 Y
port 1 e
rlabel m2 103 7 103 7 3 GND
rlabel m2 89 34 89 34 3 #10
rlabel m2 90 42 90 42 3 Y
port 1 e
rlabel m2 92 50 92 50 3 Y
port 1 e
rlabel m2 93 31 93 31 3 #10
rlabel m2c 89 50 89 50 3 Y
port 1 e
rlabel m2c 90 31 90 31 3 #10
rlabel m2 88 49 88 49 3 Y
port 1 e
rlabel m2 88 50 88 50 3 Y
port 1 e
rlabel m2 72 29 72 29 3 #10
rlabel m2 72 30 72 30 3 #10
rlabel m2 72 31 72 31 3 #10
rlabel m2 89 32 89 32 3 #10
rlabel m2 83 33 83 33 3 Y
port 1 e
rlabel m2c 69 29 69 29 3 #10
rlabel m2c 80 33 80 33 3 Y
port 1 e
rlabel m2 80 37 80 37 3 Y
port 1 e
rlabel m2 80 40 80 40 3 Y
port 1 e
rlabel m2 68 28 68 28 3 #10
rlabel m2 68 29 68 29 3 #10
rlabel m2 79 32 79 32 3 Y
port 1 e
rlabel m2 79 33 79 33 3 Y
port 1 e
rlabel m2 79 36 79 36 3 Y
port 1 e
rlabel m2 55 46 55 46 3 Y
port 1 e
rlabel m2 77 88 77 88 3 Vdd
rlabel m2 77 109 77 109 3 Vdd
rlabel m2 72 113 72 113 3 Vdd
rlabel m2 60 7 60 7 3 GND
rlabel m2 63 28 63 28 3 GND
rlabel m2 68 32 68 32 3 #10
rlabel m2c 52 46 52 46 3 Y
port 1 e
rlabel m2c 73 88 73 88 3 Vdd
rlabel m2c 73 109 73 109 3 Vdd
rlabel m2c 60 28 60 28 3 GND
rlabel m2 51 45 51 45 3 Y
port 1 e
rlabel m2 51 46 51 46 3 Y
port 1 e
rlabel m2 59 65 59 65 3 S
port 3 e
rlabel m2 72 87 72 87 3 Vdd
rlabel m2 72 88 72 88 3 Vdd
rlabel m2 72 92 72 92 3 Vdd
rlabel m2 72 109 72 109 3 Vdd
rlabel m2 59 112 59 112 3 S
port 3 e
rlabel m2 53 13 53 13 3 _S
rlabel m2 59 27 59 27 3 GND
rlabel m2 59 28 59 28 3 GND
rlabel m2 59 31 59 31 3 GND
rlabel m2 58 51 58 51 3 Y
port 1 e
rlabel m2 107 61 107 61 3 GND
rlabel m2c 55 65 55 65 3 S
port 3 e
rlabel m2c 55 112 55 112 3 S
port 3 e
rlabel m2 49 12 49 12 3 _S
rlabel m2c 50 13 50 13 3 _S
rlabel m2 52 50 52 50 3 Y
port 1 e
rlabel m2c 103 61 103 61 3 GND
rlabel m2 54 64 54 64 3 S
port 3 e
rlabel m2 54 65 54 65 3 S
port 3 e
rlabel m2 54 69 54 69 3 S
port 3 e
rlabel m2 54 112 54 112 3 S
port 3 e
rlabel m2 45 113 45 113 3 B
port 2 e
rlabel m2 42 13 42 13 3 _S
rlabel m2 42 16 42 16 3 _S
rlabel m2 42 17 42 17 3 _S
rlabel m2 51 49 51 49 3 Y
port 1 e
rlabel m2 102 60 102 60 3 GND
rlabel m2 102 61 102 61 3 GND
rlabel m2 102 65 102 65 3 GND
rlabel m2c 42 113 42 113 3 B
port 2 e
rlabel m2 45 62 45 62 3 B
port 2 e
rlabel m2 41 65 41 65 3 B
port 2 e
rlabel m2 41 113 41 113 3 B
port 2 e
rlabel m2 54 116 54 116 3 S
port 3 e
rlabel m2 44 48 44 48 3 _S
rlabel m2 52 52 52 52 3 Y
port 1 e
rlabel m2 52 53 52 53 3 Y
port 1 e
rlabel m2 52 54 52 54 3 Y
port 1 e
rlabel m2c 42 62 42 62 3 B
port 2 e
rlabel m2 24 28 24 28 3 GND
rlabel m2c 41 48 41 48 3 _S
rlabel m2 41 61 41 61 3 B
port 2 e
rlabel m2 41 62 41 62 3 B
port 2 e
rlabel m2 28 63 28 63 3 A
port 4 e
rlabel m2 28 112 28 112 3 A
port 4 e
rlabel m2 41 116 41 116 3 B
port 2 e
rlabel m2 28 29 28 29 3 GND
rlabel m2 40 47 40 47 3 _S
rlabel m2 40 48 40 48 3 _S
rlabel m2 40 51 40 51 3 _S
rlabel m2c 24 63 24 63 3 A
port 4 e
rlabel m2c 24 112 24 112 3 A
port 4 e
rlabel m2c 25 29 25 29 3 GND
rlabel m2 23 62 23 62 3 A
port 4 e
rlabel m2 23 63 23 63 3 A
port 4 e
rlabel m2 23 67 23 67 3 A
port 4 e
rlabel m2 23 112 23 112 3 A
port 4 e
rlabel m2 23 116 23 116 3 A
port 4 e
rlabel m2 14 4 14 4 3 GND
rlabel m2 14 7 14 7 3 GND
rlabel m2 14 29 14 29 3 GND
rlabel m2 14 32 14 32 3 GND
<< end >>
