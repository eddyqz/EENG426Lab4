magic
tech sky130l
timestamp 1668322234
<< ndiffusion >>
rect 8 17 13 18
rect 8 14 9 17
rect 12 14 13 17
rect 8 5 13 14
rect 15 9 20 18
rect 15 6 16 9
rect 19 6 20 9
rect 15 5 20 6
rect 22 17 27 18
rect 22 14 23 17
rect 26 14 27 17
rect 22 5 27 14
rect 34 17 39 18
rect 34 14 35 17
rect 38 14 39 17
rect 34 6 39 14
rect 41 17 48 18
rect 41 14 43 17
rect 46 14 48 17
rect 41 6 48 14
rect 50 17 55 18
rect 50 14 51 17
rect 54 14 55 17
rect 50 6 55 14
rect 62 17 67 18
rect 62 14 63 17
rect 66 14 67 17
rect 62 6 67 14
rect 69 17 76 18
rect 69 14 71 17
rect 74 14 76 17
rect 69 6 76 14
rect 78 17 83 18
rect 78 14 79 17
rect 82 14 83 17
rect 78 6 83 14
<< ndc >>
rect 9 14 12 17
rect 16 6 19 9
rect 23 14 26 17
rect 35 14 38 17
rect 43 14 46 17
rect 51 14 54 17
rect 63 14 66 17
rect 71 14 74 17
rect 79 14 82 17
<< ntransistor >>
rect 13 5 15 18
rect 20 5 22 18
rect 39 6 41 18
rect 48 6 50 18
rect 67 6 69 18
rect 76 6 78 18
<< pdiffusion >>
rect 8 29 13 42
rect 8 26 9 29
rect 12 26 13 29
rect 8 25 13 26
rect 15 41 20 42
rect 15 38 16 41
rect 19 38 20 41
rect 15 25 20 38
rect 22 29 27 42
rect 44 37 48 47
rect 22 26 23 29
rect 26 26 27 29
rect 22 25 27 26
rect 34 36 39 37
rect 34 33 35 36
rect 38 33 39 36
rect 34 25 39 33
rect 41 29 48 37
rect 41 26 43 29
rect 46 26 48 29
rect 41 25 48 26
rect 50 46 55 47
rect 50 43 51 46
rect 54 43 55 46
rect 50 25 55 43
rect 70 46 76 47
rect 70 43 71 46
rect 74 43 76 46
rect 70 37 76 43
rect 62 36 67 37
rect 62 33 63 36
rect 66 33 67 36
rect 62 25 67 33
rect 69 25 76 37
rect 78 46 83 47
rect 78 43 79 46
rect 82 43 83 46
rect 78 25 83 43
<< pdc >>
rect 9 26 12 29
rect 16 38 19 41
rect 23 26 26 29
rect 35 33 38 36
rect 43 26 46 29
rect 51 43 54 46
rect 71 43 74 46
rect 63 33 66 36
rect 79 43 82 46
<< ptransistor >>
rect 13 25 15 42
rect 20 25 22 42
rect 39 25 41 37
rect 48 25 50 47
rect 67 25 69 37
rect 76 25 78 47
<< polysilicon >>
rect 44 60 50 61
rect 44 57 45 60
rect 48 57 50 60
rect 44 55 50 57
rect 6 49 15 50
rect 6 46 7 49
rect 10 46 15 49
rect 48 47 50 55
rect 76 47 78 49
rect 6 45 15 46
rect 13 42 15 45
rect 20 42 22 44
rect 39 37 41 39
rect 67 37 69 39
rect 13 18 15 25
rect 20 18 22 25
rect 39 18 41 25
rect 48 18 50 25
rect 67 18 69 25
rect 76 22 78 25
rect 86 23 91 24
rect 86 22 87 23
rect 76 20 87 22
rect 90 20 91 23
rect 76 18 78 20
rect 86 19 91 20
rect 13 3 15 5
rect 20 -6 22 5
rect 39 3 41 6
rect 48 4 50 6
rect 67 3 69 6
rect 76 4 78 6
rect 27 2 41 3
rect 27 -1 28 2
rect 31 1 41 2
rect 62 2 69 3
rect 31 -1 32 1
rect 27 -2 32 -1
rect 62 -1 63 2
rect 66 -1 69 2
rect 62 -2 69 -1
rect 19 -7 24 -6
rect 19 -10 20 -7
rect 23 -10 24 -7
rect 19 -11 24 -10
<< pc >>
rect 45 57 48 60
rect 7 46 10 49
rect 87 20 90 23
rect 28 -1 31 2
rect 63 -1 66 2
rect 20 -10 23 -7
<< m1 >>
rect 35 70 66 73
rect 23 65 28 66
rect 23 62 24 65
rect 27 62 28 65
rect 23 61 28 62
rect 16 53 21 54
rect 16 50 17 53
rect 20 50 21 53
rect 2 49 11 50
rect 2 46 7 49
rect 10 46 11 49
rect 2 45 11 46
rect 16 49 21 50
rect 2 -23 5 45
rect 16 42 19 49
rect 15 41 20 42
rect 15 38 16 41
rect 19 38 20 41
rect 15 37 20 38
rect 24 30 27 61
rect 35 37 38 70
rect 44 65 49 66
rect 44 62 45 65
rect 48 62 49 65
rect 44 60 49 62
rect 44 57 45 60
rect 48 57 49 60
rect 44 56 49 57
rect 52 65 57 66
rect 52 62 53 65
rect 56 62 57 65
rect 52 61 57 62
rect 52 47 55 61
rect 50 46 55 47
rect 50 43 51 46
rect 54 43 55 46
rect 50 42 55 43
rect 63 37 66 70
rect 78 65 83 66
rect 78 62 79 65
rect 82 62 83 65
rect 78 61 83 62
rect 70 53 75 54
rect 70 50 71 53
rect 74 50 75 53
rect 70 46 75 50
rect 79 47 82 61
rect 70 43 71 46
rect 74 43 75 46
rect 70 42 75 43
rect 78 46 83 47
rect 78 43 79 46
rect 82 43 83 46
rect 78 42 83 43
rect 34 36 39 37
rect 34 33 35 36
rect 38 33 39 36
rect 34 32 39 33
rect 62 36 67 37
rect 62 33 63 36
rect 66 33 67 36
rect 62 32 67 33
rect 8 29 13 30
rect 8 26 9 29
rect 12 26 13 29
rect 8 25 13 26
rect 22 29 27 30
rect 22 26 23 29
rect 26 26 27 29
rect 22 25 27 26
rect 42 29 47 30
rect 42 26 43 29
rect 46 26 47 29
rect 42 25 47 26
rect 9 18 12 25
rect 23 18 26 25
rect 43 18 46 25
rect 86 23 91 24
rect 86 20 87 23
rect 90 20 91 23
rect 86 19 91 20
rect 8 17 13 18
rect 8 14 9 17
rect 12 14 13 17
rect 8 13 13 14
rect 22 17 27 18
rect 22 14 23 17
rect 26 14 27 17
rect 22 13 27 14
rect 34 17 39 18
rect 34 14 35 17
rect 38 14 39 17
rect 34 13 39 14
rect 42 17 47 18
rect 42 14 43 17
rect 46 14 47 17
rect 42 13 47 14
rect 50 17 55 18
rect 62 17 67 18
rect 50 14 51 17
rect 54 14 63 17
rect 66 14 67 17
rect 50 13 55 14
rect 62 13 67 14
rect 70 17 75 18
rect 70 14 71 17
rect 74 14 75 17
rect 70 13 75 14
rect 78 17 83 18
rect 78 14 79 17
rect 82 14 83 17
rect 78 13 83 14
rect 9 -14 12 13
rect 15 9 20 10
rect 15 6 16 9
rect 19 6 20 9
rect 15 5 20 6
rect 16 2 19 5
rect 27 2 32 3
rect 15 1 20 2
rect 15 -2 16 1
rect 19 -2 20 1
rect 27 -1 28 2
rect 31 -1 32 2
rect 27 -2 32 -1
rect 15 -3 20 -2
rect 19 -7 24 -6
rect 28 -7 31 -2
rect 35 -5 38 13
rect 19 -10 20 -7
rect 23 -10 31 -7
rect 34 -6 39 -5
rect 34 -9 35 -6
rect 38 -9 39 -6
rect 34 -10 39 -9
rect 19 -11 24 -10
rect 8 -15 13 -14
rect 8 -18 9 -15
rect 12 -18 13 -15
rect 8 -19 13 -18
rect 43 -23 46 13
rect 71 3 74 13
rect 62 2 67 3
rect 62 -1 63 2
rect 66 -1 67 2
rect 62 -2 67 -1
rect 70 2 75 3
rect 70 -1 71 2
rect 74 -1 75 2
rect 70 -2 75 -1
rect 63 -14 66 -2
rect 79 -5 82 13
rect 78 -6 83 -5
rect 78 -9 79 -6
rect 82 -9 83 -6
rect 78 -10 83 -9
rect 62 -15 67 -14
rect 62 -18 63 -15
rect 66 -18 67 -15
rect 62 -19 67 -18
rect 2 -26 46 -23
<< m2c >>
rect 24 62 27 65
rect 17 50 20 53
rect 45 62 48 65
rect 53 62 56 65
rect 79 62 82 65
rect 71 50 74 53
rect 16 -2 19 1
rect 35 -9 38 -6
rect 9 -18 12 -15
rect 71 -1 74 2
rect 79 -9 82 -6
rect 63 -18 66 -15
<< m2 >>
rect 23 65 28 66
rect 44 65 49 66
rect 23 62 24 65
rect 27 62 45 65
rect 48 62 49 65
rect 23 61 28 62
rect 44 61 49 62
rect 52 65 57 66
rect 78 65 83 66
rect 52 62 53 65
rect 56 62 79 65
rect 82 62 83 65
rect 52 61 57 62
rect 78 61 83 62
rect 16 53 21 54
rect 70 53 75 54
rect 16 50 17 53
rect 20 50 71 53
rect 74 50 75 53
rect 16 49 21 50
rect 70 49 75 50
rect 70 2 75 3
rect 15 1 71 2
rect 15 -2 16 1
rect 19 -1 71 1
rect 74 -1 75 2
rect 19 -2 20 -1
rect 70 -2 75 -1
rect 15 -3 20 -2
rect 34 -6 39 -5
rect 78 -6 83 -5
rect 34 -9 35 -6
rect 38 -9 79 -6
rect 82 -9 83 -6
rect 34 -10 39 -9
rect 78 -10 83 -9
rect 8 -15 13 -14
rect 62 -15 67 -14
rect 8 -18 9 -15
rect 12 -18 63 -15
rect 66 -18 67 -15
rect 8 -19 13 -18
rect 62 -19 67 -18
<< labels >>
rlabel ndiffusion 51 7 51 7 3 #10
rlabel ntransistor 49 17 49 17 3 _clk
rlabel ndiffusion 42 7 42 7 3 _q
rlabel ntransistor 40 17 40 17 3 CLK
rlabel ndiffusion 35 7 35 7 3 #5
rlabel ndiffusion 79 7 79 7 3 #5
rlabel ntransistor 77 17 77 17 3 D
rlabel ndiffusion 70 7 70 7 3 GND
rlabel ntransistor 68 17 68 17 3 Q
rlabel ndiffusion 63 7 63 7 3 #10
rlabel ptransistor 49 26 49 26 3 _clk
rlabel ptransistor 40 26 40 26 3 CLK
rlabel ptransistor 77 26 77 26 3 D
rlabel ptransistor 68 26 68 26 3 Q
rlabel ndiffusion 23 6 23 6 3 _clk
rlabel ntransistor 21 16 21 16 3 CLK
rlabel ndiffusion 16 6 16 6 3 GND
rlabel ntransistor 14 16 14 16 3 _q
rlabel ndiffusion 9 6 9 6 3 Q
rlabel ptransistor 21 26 21 26 3 CLK
rlabel ptransistor 14 26 14 26 3 _q
rlabel m1 44 71 44 71 5 #8
rlabel m2 43 51 43 51 1 Vdd
rlabel m2 72 64 72 64 1 #7
rlabel m2 53 1 53 1 1 GND
rlabel m2 56 -7 56 -7 1 #5
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 88 52
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
