magic
tech sky130l
timestamp 1668327865
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 12 19 15
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 28 13 53
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 23 20 53
rect 22 28 27 53
rect 22 25 23 28
rect 26 25 27 28
rect 22 23 27 25
<< pdc >>
rect 9 25 12 28
rect 23 25 26 28
<< ptransistor >>
rect 13 23 15 53
rect 20 23 22 53
<< polysilicon >>
rect 10 61 15 62
rect 10 58 11 61
rect 14 58 15 61
rect 10 57 15 58
rect 13 53 15 57
rect 20 61 25 62
rect 20 58 21 61
rect 24 58 25 61
rect 20 57 25 58
rect 20 53 22 57
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 11 58 14 61
rect 21 58 24 61
<< m1 >>
rect 10 61 15 62
rect 10 58 11 61
rect 14 58 15 61
rect 10 57 15 58
rect 20 61 25 62
rect 20 58 21 61
rect 24 58 25 61
rect 20 57 25 58
rect 3 28 13 29
rect 3 25 4 28
rect 7 25 9 28
rect 12 25 13 28
rect 3 24 13 25
rect 23 28 26 29
rect 23 21 26 25
rect 16 18 26 21
rect 16 15 19 18
rect 16 11 19 12
rect 9 10 12 11
rect 9 4 12 7
rect 23 10 26 11
rect 23 4 26 7
rect 8 3 13 4
rect 8 0 9 3
rect 12 0 13 3
rect 8 -1 13 0
rect 22 3 27 4
rect 22 0 23 3
rect 26 0 27 3
rect 22 -1 27 0
<< m2c >>
rect 4 25 7 28
rect 9 0 12 3
rect 23 0 26 3
<< m2 >>
rect 1 28 8 29
rect 1 25 4 28
rect 7 25 8 28
rect 1 24 8 25
rect 8 3 13 4
rect 22 3 27 4
rect 8 0 9 3
rect 12 0 23 3
rect 26 0 27 3
rect 8 -1 13 0
rect 22 -1 27 0
<< labels >>
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 17 21 17 3 B
rlabel polysilicon 21 22 21 22 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 18 19 18 19 1 Y
rlabel m2 17 1 17 1 1 GND
rlabel m2 2 27 2 27 3 Vdd
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 40 64
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
