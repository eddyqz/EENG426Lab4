magic
tech sky130l
timestamp 1668469005
<< checkpaint >>
rect -24 92 108 100
rect -24 84 109 92
rect -30 23 109 84
rect -30 17 108 23
rect -30 -14 104 17
rect -24 -18 104 -14
rect -24 -24 103 -18
rect -24 -25 100 -24
rect -24 -28 64 -25
rect -24 -29 48 -28
rect -24 -30 43 -29
<< ndiffusion >>
rect 8 21 13 24
rect 8 18 9 21
rect 12 18 13 21
rect 8 14 13 18
rect 15 14 20 24
rect 22 20 27 24
rect 22 17 23 20
rect 26 17 27 20
rect 22 14 27 17
rect 34 20 39 24
rect 34 17 35 20
rect 38 17 39 20
rect 34 14 39 17
rect 41 18 46 24
rect 41 15 42 18
rect 45 15 46 18
rect 41 14 46 15
rect 48 22 53 24
rect 48 19 49 22
rect 52 19 53 22
rect 48 14 53 19
rect 60 21 65 24
rect 60 18 61 21
rect 64 18 65 21
rect 60 14 65 18
rect 67 21 72 24
rect 67 18 68 21
rect 71 18 72 21
rect 67 14 72 18
<< ndc >>
rect 9 18 12 21
rect 23 17 26 20
rect 35 17 38 20
rect 42 15 45 18
rect 49 19 52 22
rect 61 18 64 21
rect 68 18 71 21
<< ntransistor >>
rect 13 14 15 24
rect 20 14 22 24
rect 39 14 41 24
rect 46 14 48 24
rect 65 14 67 24
<< pdiffusion >>
rect 8 46 13 51
rect 8 43 9 46
rect 12 43 13 46
rect 8 31 13 43
rect 15 46 19 51
rect 15 38 20 46
rect 15 35 16 38
rect 19 35 20 38
rect 15 31 20 35
rect 22 37 27 46
rect 60 46 65 51
rect 60 43 61 46
rect 64 43 65 46
rect 22 34 23 37
rect 26 34 27 37
rect 22 31 27 34
rect 34 37 39 41
rect 34 34 35 37
rect 38 34 39 37
rect 34 31 39 34
rect 41 31 46 41
rect 48 38 53 41
rect 48 35 49 38
rect 52 35 53 38
rect 48 31 53 35
rect 60 31 65 43
rect 67 36 72 51
rect 67 33 68 36
rect 71 33 72 36
rect 67 31 72 33
<< pdc >>
rect 9 43 12 46
rect 16 35 19 38
rect 61 43 64 46
rect 23 34 26 37
rect 35 34 38 37
rect 49 35 52 38
rect 68 33 71 36
<< ptransistor >>
rect 13 31 15 51
rect 20 31 22 46
rect 39 31 41 41
rect 46 31 48 41
rect 65 31 67 51
<< polysilicon >>
rect 16 66 21 67
rect 16 63 17 66
rect 20 64 21 66
rect 20 63 22 64
rect 46 63 48 64
rect 16 62 22 63
rect 12 58 17 59
rect 12 55 13 58
rect 16 55 17 58
rect 12 54 17 55
rect 13 51 15 54
rect 20 50 22 62
rect 43 62 49 63
rect 43 58 44 62
rect 48 58 49 62
rect 43 57 49 58
rect 20 48 41 50
rect 20 46 22 48
rect 39 41 41 48
rect 46 41 48 57
rect 65 51 67 53
rect 13 24 15 31
rect 20 24 22 31
rect 39 24 41 31
rect 46 24 48 31
rect 65 24 67 31
rect 13 12 15 14
rect 20 12 22 14
rect 39 12 41 14
rect 46 12 48 14
rect 65 12 67 14
rect 63 11 68 12
rect 63 8 64 11
rect 67 8 68 11
rect 63 7 68 8
<< pc >>
rect 17 63 20 66
rect 13 55 16 58
rect 44 58 48 62
rect 64 8 67 11
<< m1 >>
rect 8 67 12 68
rect 8 66 21 67
rect 8 64 17 66
rect 16 63 17 64
rect 20 63 21 66
rect 16 62 21 63
rect 24 64 28 68
rect 12 58 17 59
rect 24 58 27 64
rect 12 55 13 58
rect 16 55 27 58
rect 40 63 44 68
rect 52 67 60 68
rect 52 64 53 67
rect 56 64 60 67
rect 72 64 76 68
rect 52 63 57 64
rect 40 62 49 63
rect 40 58 44 62
rect 48 58 49 62
rect 40 57 49 58
rect 73 59 76 64
rect 73 52 76 56
rect 2 49 76 52
rect 2 21 5 49
rect 8 43 9 46
rect 12 43 61 46
rect 64 43 65 46
rect 16 38 19 39
rect 49 38 52 39
rect 35 37 38 38
rect 16 34 19 35
rect 22 34 23 37
rect 26 34 32 37
rect 2 18 9 21
rect 12 18 13 21
rect 23 20 26 21
rect 23 16 26 17
rect 29 20 32 34
rect 49 34 52 35
rect 68 36 71 37
rect 35 33 38 34
rect 68 32 71 33
rect 49 26 71 29
rect 49 22 52 26
rect 29 17 35 20
rect 38 17 39 20
rect 42 18 45 19
rect 49 18 52 19
rect 61 21 64 22
rect 29 11 32 17
rect 61 17 64 18
rect 68 21 71 26
rect 68 17 71 18
rect 42 14 45 15
rect 63 11 68 12
rect 29 8 64 11
rect 67 8 68 11
rect 63 7 68 8
rect 8 4 12 7
rect 15 4 16 7
rect 8 2 11 4
<< m2c >>
rect 53 64 56 67
rect 73 56 76 59
rect 16 35 19 38
rect 23 17 26 20
rect 35 34 38 37
rect 49 35 52 38
rect 68 33 71 36
rect 61 18 64 21
rect 42 15 45 18
rect 12 4 15 7
<< m2 >>
rect 49 67 57 68
rect 49 64 53 67
rect 56 64 57 67
rect 49 63 57 64
rect 49 62 52 63
rect 16 59 52 62
rect 16 39 19 59
rect 49 39 52 59
rect 72 59 77 60
rect 72 58 73 59
rect 55 56 73 58
rect 76 56 77 59
rect 15 38 20 39
rect 48 38 53 39
rect 15 35 16 38
rect 19 35 20 38
rect 15 34 20 35
rect 29 37 39 38
rect 29 34 35 37
rect 38 34 39 37
rect 48 35 49 38
rect 52 35 53 38
rect 48 34 53 35
rect 29 33 39 34
rect 22 20 27 21
rect 29 20 32 33
rect 22 17 23 20
rect 26 17 32 20
rect 22 16 27 17
rect 29 11 32 17
rect 41 18 46 19
rect 41 15 42 18
rect 45 16 46 18
rect 55 16 57 56
rect 72 55 77 56
rect 67 36 72 37
rect 67 33 68 36
rect 71 33 72 36
rect 67 32 72 33
rect 60 21 65 22
rect 60 18 61 21
rect 64 18 65 21
rect 60 17 65 18
rect 45 15 57 16
rect 41 14 57 15
rect 61 11 64 17
rect 68 11 71 32
rect 29 8 71 11
rect 11 7 16 8
rect 29 7 32 8
rect 11 4 12 7
rect 15 4 32 7
rect 11 3 16 4
<< labels >>
rlabel ndiffusion 72 19 72 19 3 #10
rlabel ndiffusion 68 15 68 15 3 #10
rlabel ndiffusion 68 19 68 19 3 #10
rlabel ndiffusion 68 22 68 22 3 #10
rlabel pdiffusion 68 32 68 32 3 _q
rlabel ntransistor 66 15 66 15 3 _clk
rlabel polysilicon 66 25 66 25 3 _clk
rlabel ptransistor 66 32 66 32 3 _clk
rlabel polysilicon 66 52 66 52 3 _clk
rlabel ndiffusion 61 15 61 15 3 _q
rlabel ndiffusion 53 20 53 20 3 #10
rlabel pdiffusion 61 32 61 32 3 #7
rlabel pdiffusion 61 44 61 44 3 #7
rlabel pdiffusion 61 47 61 47 3 #7
rlabel ndiffusion 49 15 49 15 3 #10
rlabel ndiffusion 49 20 49 20 3 #10
rlabel ndiffusion 49 23 49 23 3 #10
rlabel pdiffusion 49 32 49 32 3 Vdd
rlabel polysilicon 47 42 47 42 3 q
rlabel polysilicon 47 64 47 64 3 q
rlabel polysilicon 66 13 66 13 3 _clk
rlabel ntransistor 47 15 47 15 3 q
rlabel polysilicon 47 25 47 25 3 q
rlabel ptransistor 47 32 47 32 3 q
rlabel polysilicon 44 58 44 58 3 q
rlabel polysilicon 44 59 44 59 3 q
rlabel polysilicon 44 63 44 63 3 q
rlabel ndiffusion 35 18 35 18 3 _clk
rlabel polysilicon 47 13 47 13 3 q
rlabel ntransistor 40 15 40 15 3 CLK
rlabel polysilicon 40 25 40 25 3 CLK
rlabel ptransistor 40 32 40 32 3 CLK
rlabel polysilicon 40 42 40 42 3 CLK
rlabel ndiffusion 35 15 35 15 3 _clk
rlabel ndiffusion 35 21 35 21 3 _clk
rlabel pdiffusion 35 32 35 32 3 _q
rlabel pdiffusion 35 35 35 35 3 _q
rlabel pdiffusion 35 38 35 38 3 _q
rlabel polysilicon 21 65 21 65 3 CLK
rlabel polysilicon 40 13 40 13 3 CLK
rlabel ndiffusion 23 15 23 15 3 _q
rlabel pdiffusion 23 32 23 32 3 _clk
rlabel pdiffusion 23 38 23 38 3 _clk
rlabel polysilicon 21 47 21 47 3 CLK
rlabel polysilicon 21 49 21 49 3 CLK
rlabel polysilicon 21 51 21 51 3 CLK
rlabel polysilicon 17 67 17 67 3 CLK
rlabel polysilicon 21 13 21 13 3 CLK
rlabel ntransistor 21 15 21 15 3 CLK
rlabel polysilicon 21 25 21 25 3 CLK
rlabel ptransistor 21 32 21 32 3 CLK
rlabel polysilicon 64 9 64 9 3 _clk
rlabel pdiffusion 16 32 16 32 3 Vdd
rlabel pdiffusion 16 47 16 47 3 Vdd
rlabel polysilicon 14 52 14 52 3 D
rlabel polysilicon 14 13 14 13 3 D
rlabel ntransistor 14 15 14 15 3 D
rlabel polysilicon 14 25 14 25 3 D
rlabel ptransistor 14 32 14 32 3 D
rlabel polysilicon 13 55 13 55 3 D
rlabel ndiffusion 9 15 9 15 3 GND
rlabel ndiffusion 9 19 9 19 3 GND
rlabel ndiffusion 9 22 9 22 3 GND
rlabel pdiffusion 9 32 9 32 3 #7
rlabel pdiffusion 9 47 9 47 3 #7
rlabel m1 74 53 74 53 3 GND
rlabel m1 74 60 74 60 3 GND
rlabel m1 73 65 73 65 3 GND
rlabel ndc 69 19 69 19 3 #10
rlabel m1 69 22 69 22 3 #10
rlabel m1 69 33 69 33 3 _q
port 1 e
rlabel m1 69 37 69 37 3 _q
port 1 e
rlabel m1 62 22 62 22 3 _q
port 1 e
rlabel m1 53 64 53 64 3 Vdd
rlabel m1 53 65 53 65 3 Vdd
rlabel m1 53 68 53 68 3 Vdd
rlabel m1 49 59 49 59 3 q
port 2 e
rlabel m1 50 19 50 19 3 #10
rlabel ndc 50 20 50 20 3 #10
rlabel m1 50 23 50 23 3 #10
rlabel m1 50 27 50 27 3 #10
rlabel m1 50 35 50 35 3 Vdd
rlabel m1 50 39 50 39 3 Vdd
rlabel pc 45 59 45 59 3 q
port 2 e
rlabel m1 41 58 41 58 3 q
port 2 e
rlabel m1 41 59 41 59 3 q
port 2 e
rlabel m1 41 63 41 63 3 q
port 2 e
rlabel m1 41 64 41 64 3 q
port 2 e
rlabel m1 43 19 43 19 3 GND
rlabel m1 69 18 69 18 3 #10
rlabel m1 36 38 36 38 3 _q
port 1 e
rlabel m1 39 18 39 18 3 _clk
rlabel m1 36 34 36 34 3 _q
port 1 e
rlabel m1 62 18 62 18 3 _q
port 1 e
rlabel ndc 36 18 36 18 3 _clk
rlabel m1 27 35 27 35 3 _clk
rlabel m1 64 12 64 12 3 _clk
rlabel m1 30 18 30 18 3 _clk
rlabel m1 30 21 30 21 3 _clk
rlabel pdc 24 35 24 35 3 _clk
rlabel m1 25 59 25 59 3 D
port 3 e
rlabel m1 25 65 25 65 3 D
port 3 e
rlabel m1 21 64 21 64 3 CLK
port 4 e
rlabel m1 64 8 64 8 3 _clk
rlabel m1 68 9 68 9 3 _clk
rlabel m1 43 15 43 15 3 GND
rlabel m1 23 35 23 35 3 _clk
rlabel m1 65 44 65 44 3 #7
rlabel pc 18 64 18 64 3 CLK
port 4 e
rlabel pc 65 9 65 9 3 _clk
rlabel m1 24 17 24 17 3 _q
port 1 e
rlabel m1 24 21 24 21 3 _q
port 1 e
rlabel pdc 62 44 62 44 3 #7
rlabel m1 17 56 17 56 3 D
port 3 e
rlabel m1 17 63 17 63 3 CLK
port 4 e
rlabel m1 17 64 17 64 3 CLK
port 4 e
rlabel m1 30 9 30 9 3 _clk
rlabel m1 30 12 30 12 3 _clk
rlabel m1 17 35 17 35 3 Vdd
rlabel m1 17 39 17 39 3 Vdd
rlabel m1 13 44 13 44 3 #7
rlabel pc 14 56 14 56 3 D
port 3 e
rlabel pdc 10 44 10 44 3 #7
rlabel m1 13 56 13 56 3 D
port 3 e
rlabel m1 13 59 13 59 3 D
port 3 e
rlabel m1 13 19 13 19 3 GND
rlabel m1 9 44 9 44 3 #7
rlabel m1 9 3 9 3 3 _q
port 1 e
rlabel m1 9 5 9 5 3 _q
port 1 e
rlabel ndc 10 19 10 19 3 GND
rlabel m1 9 65 9 65 3 CLK
port 4 e
rlabel m1 9 67 9 67 3 CLK
port 4 e
rlabel m1 9 68 9 68 3 CLK
port 4 e
rlabel m1 3 19 3 19 3 GND
rlabel m1 3 22 3 22 3 GND
rlabel m1 3 50 3 50 3 GND
rlabel m2 73 56 73 56 3 GND
rlabel m2 72 34 72 34 3 _q
port 1 e
rlabel m2c 69 34 69 34 3 _q
port 1 e
rlabel m2 73 59 73 59 3 GND
rlabel m2 73 60 73 60 3 GND
rlabel m2 65 19 65 19 3 _q
port 1 e
rlabel m2 68 33 68 33 3 _q
port 1 e
rlabel m2 68 34 68 34 3 _q
port 1 e
rlabel m2 68 37 68 37 3 _q
port 1 e
rlabel m2c 62 19 62 19 3 _q
port 1 e
rlabel m2 61 18 61 18 3 _q
port 1 e
rlabel m2 61 19 61 19 3 _q
port 1 e
rlabel m2 61 22 61 22 3 _q
port 1 e
rlabel m2 77 57 77 57 3 GND
rlabel m2 69 12 69 12 3 _q
port 1 e
rlabel m2c 74 57 74 57 3 GND
rlabel m2 56 17 56 17 3 GND
rlabel m2 56 57 56 57 3 GND
rlabel m2 62 12 62 12 3 _q
port 1 e
rlabel m2 53 36 53 36 3 Vdd
rlabel m2c 50 36 50 36 3 Vdd
rlabel m2 50 40 50 40 3 Vdd
rlabel m2 57 65 57 65 3 Vdd
rlabel m2 46 16 46 16 3 GND
rlabel m2 46 17 46 17 3 GND
rlabel m2 49 35 49 35 3 Vdd
rlabel m2 49 36 49 36 3 Vdd
rlabel m2 49 39 49 39 3 Vdd
rlabel m2c 54 65 54 65 3 Vdd
rlabel m2c 43 16 43 16 3 GND
rlabel m2 42 19 42 19 3 GND
rlabel m2 50 63 50 63 3 Vdd
rlabel m2 50 64 50 64 3 Vdd
rlabel m2 50 65 50 65 3 Vdd
rlabel m2 50 68 50 68 3 Vdd
rlabel m2 42 15 42 15 3 GND
rlabel m2 42 16 42 16 3 GND
rlabel m2 39 35 39 35 3 _q
port 1 e
rlabel m2 30 38 30 38 3 _q
port 1 e
rlabel m2c 36 35 36 35 3 _q
port 1 e
rlabel m2 30 8 30 8 3 _q
port 1 e
rlabel m2 30 9 30 9 3 _q
rlabel m2 30 12 30 12 3 _q
rlabel m2 27 18 27 18 3 _q
port 1 e
rlabel m2 30 21 30 21 3 _q
rlabel m2 30 34 30 34 3 _q
port 1 e
rlabel m2 30 35 30 35 3 _q
port 1 e
rlabel m2 20 36 20 36 3 Vdd
rlabel m2c 24 18 24 18 3 _q
port 1 e
rlabel m2c 17 36 17 36 3 Vdd
rlabel m2 17 40 17 40 3 Vdd
rlabel m2 17 60 17 60 3 Vdd
rlabel m2 16 5 16 5 3 _q
port 1 e
rlabel m2 23 17 23 17 3 _q
port 1 e
rlabel m2 23 18 23 18 3 _q
port 1 e
rlabel m2 23 21 23 21 3 _q
port 1 e
rlabel m2 16 35 16 35 3 Vdd
rlabel m2 16 36 16 36 3 Vdd
rlabel m2 16 39 16 39 3 Vdd
rlabel m2c 13 5 13 5 3 _q
port 1 e
rlabel m2 12 4 12 4 3 _q
port 1 e
rlabel m2 12 5 12 5 3 _q
port 1 e
rlabel m2 12 8 12 8 3 _q
port 1 e
<< end >>
