VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.600000 BY 0.300000 ;
END CoreSite

LAYER li1
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.056250 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.225000 ;
   PITCH 0.600000 0.600000 ;
END li1

LAYER mcon
    TYPE CUT ;
    SPACING 0.225000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END mcon

LAYER met1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.150000 ;
   AREA 0.084375 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met1

LAYER v1
    TYPE CUT ;
    SPACING 0.075000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.075000 ;
END v1

LAYER met2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.150000 ;
   AREA 0.073125 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met2

LAYER v2
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v2

LAYER met3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met3

LAYER v3
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.450000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v3

LAYER met4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met4

LAYER v4
    TYPE CUT ;
    SPACING 0.450000 ;
    WIDTH 1.200000 ;
    ENCLOSURE ABOVE 0.150000 0.150000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END v4

LAYER met5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.650000 ;
   AREA 4.005000 ;
   WIDTH 1.650000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 1.650000 ;
   PITCH 3.300000 3.300000 ;
END met5

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA mcon_C DEFAULT
   LAYER li1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER mcon ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END mcon_C

VIA v1_C DEFAULT
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER met2 ;
     RECT -0.225000 -0.150000 0.225000 0.150000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_C

VIA v3_Ch
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Ch

VIA v3_Cv
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER met4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER met5 ;
     RECT -0.750000 -0.750000 0.750000 0.750000 ;
END v4_C

MACRO _0_0std_0_0cells_0_0MUX2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0MUX2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 8.400000 BY 9.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li1 ;
        RECT 1.650000 8.625000 2.100000 8.700000 ;
        RECT 1.650000 8.325000 1.725000 8.625000 ;
        RECT 1.650000 8.250000 2.100000 8.325000 ;
        RECT 1.650000 4.950000 2.100000 5.025000 ;
        RECT 1.650000 4.650000 1.725000 4.950000 ;
        RECT 1.650000 4.575000 2.100000 4.650000 ;
        RECT 1.725000 8.325000 2.025000 8.625000 ;
        RECT 1.725000 4.650000 2.025000 4.950000 ;
        RECT 2.025000 8.325000 2.100000 8.625000 ;
        RECT 2.025000 4.650000 2.100000 4.950000 ;
        RECT 1.800000 4.500000 2.100000 4.575000 ;
        LAYER mcon ;
        RECT 1.725000 8.325000 2.025000 8.625000 ;
        RECT 1.725000 4.650000 2.025000 4.950000 ;
        LAYER met1 ;
        RECT 1.650000 8.625000 2.100000 8.700000 ;
        RECT 1.650000 8.325000 1.725000 8.625000 ;
        RECT 1.650000 4.950000 2.100000 8.325000 ;
        RECT 1.650000 4.650000 1.725000 4.950000 ;
        RECT 1.650000 4.575000 2.100000 4.650000 ;
        RECT 1.725000 8.325000 2.025000 8.625000 ;
        RECT 1.725000 4.650000 2.025000 4.950000 ;
        RECT 2.025000 8.325000 2.100000 8.625000 ;
        RECT 2.025000 4.650000 2.100000 4.950000 ;
        END
        ANTENNAGATEAREA 0.281250 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li1 ;
        RECT 3.000000 6.075000 4.650000 6.375000 ;
        RECT 3.000000 4.800000 3.300000 6.075000 ;
        RECT 3.000000 4.575000 3.075000 4.800000 ;
        RECT 3.000000 4.500000 3.300000 4.575000 ;
        RECT 4.650000 6.075000 4.950000 6.375000 ;
        RECT 3.075000 4.575000 3.300000 4.800000 ;
        RECT 3.000000 8.625000 3.375000 8.700000 ;
        RECT 3.000000 8.400000 3.075000 8.625000 ;
        RECT 3.000000 8.325000 3.375000 8.400000 ;
        RECT 4.950000 6.075000 5.025000 6.375000 ;
        RECT 3.075000 8.400000 3.300000 8.625000 ;
        RECT 3.300000 8.400000 3.375000 8.625000 ;
        RECT 4.575000 6.375000 5.025000 6.450000 ;
        RECT 4.575000 6.000000 5.025000 6.075000 ;
        LAYER mcon ;
        RECT 3.075000 8.400000 3.300000 8.625000 ;
        RECT 3.075000 4.575000 3.300000 4.800000 ;
        LAYER met1 ;
        RECT 3.000000 8.625000 3.375000 8.700000 ;
        RECT 3.000000 8.400000 3.075000 8.625000 ;
        RECT 3.000000 4.800000 3.375000 8.400000 ;
        RECT 3.000000 4.575000 3.075000 4.800000 ;
        RECT 3.000000 4.500000 3.375000 4.575000 ;
        RECT 3.075000 8.400000 3.300000 8.625000 ;
        RECT 3.075000 4.575000 3.300000 4.800000 ;
        RECT 3.300000 8.400000 3.375000 8.625000 ;
        RECT 3.300000 4.575000 3.375000 4.800000 ;
        END
        ANTENNAGATEAREA 0.281250 ;
    END B
    PIN S
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li1 ;
        RECT 3.975000 5.100000 4.425000 5.175000 ;
        RECT 3.975000 4.800000 4.050000 5.100000 ;
        RECT 3.975000 4.725000 4.500000 4.800000 ;
        RECT 4.200000 4.500000 4.500000 4.725000 ;
        RECT 4.050000 4.800000 4.350000 5.100000 ;
        RECT 3.975000 8.625000 4.425000 8.700000 ;
        RECT 3.975000 8.325000 4.050000 8.625000 ;
        RECT 3.975000 8.250000 4.425000 8.325000 ;
        RECT 4.350000 4.800000 4.425000 5.100000 ;
        RECT 4.050000 8.325000 4.350000 8.625000 ;
        RECT 4.350000 8.325000 4.425000 8.625000 ;
        LAYER mcon ;
        RECT 4.050000 8.325000 4.350000 8.625000 ;
        RECT 4.050000 4.800000 4.350000 5.100000 ;
        LAYER met1 ;
        RECT 3.975000 8.625000 4.425000 8.700000 ;
        RECT 3.975000 8.325000 4.050000 8.625000 ;
        RECT 3.975000 5.100000 4.425000 8.325000 ;
        RECT 3.975000 4.800000 4.050000 5.100000 ;
        RECT 3.975000 4.725000 4.425000 4.800000 ;
        RECT 4.050000 8.325000 4.350000 8.625000 ;
        RECT 4.050000 4.800000 4.350000 5.100000 ;
        RECT 4.350000 8.325000 4.425000 8.625000 ;
        RECT 4.350000 4.800000 4.425000 5.100000 ;
        END
        ANTENNAGATEAREA 0.438750 ;
    END S
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li1 ;
        RECT 0.675000 1.050000 3.225000 1.275000 ;
        RECT 0.675000 0.975000 1.875000 1.050000 ;
        RECT 2.850000 2.025000 3.225000 2.100000 ;
        RECT 2.850000 2.325000 3.300000 2.400000 ;
        RECT 2.850000 2.100000 2.925000 2.325000 ;
        RECT 2.925000 2.100000 3.150000 2.325000 ;
        RECT 3.000000 1.275000 3.225000 2.025000 ;
        RECT 3.150000 2.175000 3.300000 2.325000 ;
        RECT 3.150000 2.100000 3.225000 2.175000 ;
        RECT 3.075000 2.850000 3.675000 3.000000 ;
        RECT 3.075000 2.775000 3.525000 2.850000 ;
        RECT 3.075000 2.400000 3.300000 2.775000 ;
        RECT 3.300000 3.000000 3.675000 3.075000 ;
        RECT 3.450000 3.375000 3.825000 3.600000 ;
        RECT 3.450000 3.300000 4.125000 3.375000 ;
        RECT 3.450000 3.075000 3.675000 3.300000 ;
        RECT 3.825000 3.375000 4.050000 3.600000 ;
        RECT 3.750000 3.600000 4.125000 3.675000 ;
        RECT 4.050000 3.375000 4.125000 3.600000 ;
        RECT 5.850000 2.625000 6.225000 2.700000 ;
        RECT 5.850000 2.400000 5.925000 2.625000 ;
        RECT 5.850000 2.325000 6.225000 2.400000 ;
        RECT 5.925000 2.400000 6.150000 2.625000 ;
        RECT 6.150000 2.400000 6.225000 2.625000 ;
        RECT 6.525000 3.900000 6.900000 3.975000 ;
        RECT 6.525000 3.675000 6.600000 3.900000 ;
        RECT 6.525000 3.600000 6.900000 3.675000 ;
        RECT 6.600000 3.675000 6.825000 3.900000 ;
        RECT 6.825000 3.675000 6.900000 3.900000 ;
        LAYER mcon ;
        RECT 3.825000 3.375000 4.050000 3.600000 ;
        RECT 5.925000 2.400000 6.150000 2.625000 ;
        RECT 6.600000 3.675000 6.825000 3.900000 ;
        LAYER met1 ;
        RECT 3.750000 3.600000 4.125000 3.675000 ;
        RECT 3.750000 3.375000 3.825000 3.600000 ;
        RECT 3.750000 3.300000 4.125000 3.375000 ;
        RECT 3.825000 3.975000 4.275000 4.050000 ;
        RECT 3.825000 3.900000 6.900000 3.975000 ;
        RECT 3.825000 3.825000 6.600000 3.900000 ;
        RECT 3.825000 3.675000 4.050000 3.825000 ;
        RECT 3.825000 3.375000 4.050000 3.600000 ;
        RECT 4.050000 3.375000 4.125000 3.600000 ;
        RECT 4.275000 3.750000 6.600000 3.825000 ;
        RECT 5.850000 2.625000 6.225000 2.700000 ;
        RECT 5.850000 2.400000 5.925000 2.625000 ;
        RECT 5.850000 2.325000 6.225000 2.400000 ;
        RECT 5.925000 2.925000 6.825000 3.075000 ;
        RECT 5.925000 2.700000 6.150000 2.925000 ;
        RECT 5.925000 2.400000 6.150000 2.625000 ;
        RECT 6.150000 2.400000 6.225000 2.625000 ;
        RECT 6.525000 3.675000 6.600000 3.750000 ;
        RECT 6.525000 3.600000 6.900000 3.675000 ;
        RECT 6.600000 3.675000 6.825000 3.900000 ;
        RECT 6.825000 3.675000 6.900000 3.900000 ;
        RECT 6.675000 3.075000 6.825000 3.600000 ;
        END
        ANTENNADIFFAREA 1.575000 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li1 ;
        RECT 2.400000 3.750000 2.625000 6.825000 ;
        RECT 2.400000 3.525000 2.625000 3.750000 ;
        RECT 2.400000 3.450000 2.625000 3.525000 ;
        RECT 2.400000 6.825000 5.700000 7.050000 ;
        RECT 4.950000 4.200000 5.325000 4.275000 ;
        RECT 4.950000 3.975000 5.025000 4.200000 ;
        RECT 4.950000 3.900000 5.325000 3.975000 ;
        RECT 5.025000 3.975000 5.250000 4.200000 ;
        RECT 5.100000 4.500000 5.700000 4.800000 ;
        RECT 5.100000 4.275000 5.325000 4.500000 ;
        RECT 5.250000 3.975000 5.325000 4.200000 ;
        RECT 5.400000 6.525000 5.700000 6.825000 ;
        RECT 5.400000 6.150000 5.700000 6.525000 ;
        RECT 5.475000 4.800000 5.700000 6.150000 ;
        RECT 5.325000 8.400000 5.775000 8.475000 ;
        RECT 5.325000 8.100000 5.400000 8.400000 ;
        RECT 5.325000 8.025000 5.775000 8.100000 ;
        RECT 5.400000 8.100000 5.700000 8.400000 ;
        RECT 5.700000 8.100000 5.775000 8.400000 ;
        LAYER mcon ;
        RECT 5.400000 8.100000 5.700000 8.400000 ;
        RECT 5.400000 6.525000 5.700000 6.825000 ;
        LAYER met1 ;
        RECT 5.325000 8.400000 5.775000 8.475000 ;
        RECT 5.325000 8.100000 5.400000 8.400000 ;
        RECT 5.325000 6.825000 5.775000 8.100000 ;
        RECT 5.325000 6.525000 5.400000 6.825000 ;
        RECT 5.325000 6.450000 5.775000 6.525000 ;
        RECT 5.400000 8.100000 5.700000 8.400000 ;
        RECT 5.400000 6.525000 5.700000 6.825000 ;
        RECT 5.700000 8.100000 5.775000 8.400000 ;
        RECT 5.700000 6.525000 5.775000 6.825000 ;
        END
        ANTENNADIFFAREA 0.804375 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li1 ;
        RECT 1.725000 2.325000 2.100000 2.400000 ;
        RECT 1.725000 2.100000 1.800000 2.325000 ;
        RECT 1.725000 2.025000 2.100000 2.100000 ;
        RECT 1.800000 2.100000 2.025000 2.325000 ;
        RECT 2.025000 2.100000 2.100000 2.325000 ;
        RECT 4.350000 2.250000 4.725000 2.325000 ;
        RECT 4.350000 2.025000 4.425000 2.250000 ;
        RECT 4.350000 1.950000 4.725000 2.025000 ;
        RECT 4.425000 2.025000 4.650000 2.250000 ;
        RECT 4.650000 2.025000 4.725000 2.250000 ;
        RECT 7.575000 4.800000 8.025000 4.875000 ;
        RECT 6.600000 4.500000 7.650000 4.800000 ;
        RECT 7.650000 4.500000 7.950000 4.800000 ;
        RECT 7.950000 4.500000 8.025000 4.800000 ;
        RECT 7.575000 4.425000 8.025000 4.500000 ;
        LAYER mcon ;
        RECT 1.800000 2.100000 2.025000 2.325000 ;
        RECT 4.425000 2.025000 4.650000 2.250000 ;
        RECT 7.650000 4.500000 7.950000 4.800000 ;
        LAYER met1 ;
        RECT 0.975000 2.325000 2.100000 2.400000 ;
        RECT 0.975000 2.100000 1.800000 2.325000 ;
        RECT 0.975000 0.450000 1.275000 2.100000 ;
        RECT 0.975000 0.225000 7.950000 0.450000 ;
        RECT 1.800000 2.100000 2.025000 2.325000 ;
        RECT 2.025000 2.100000 2.100000 2.325000 ;
        RECT 1.725000 2.025000 2.100000 2.100000 ;
        RECT 4.350000 2.250000 4.725000 2.325000 ;
        RECT 4.350000 2.025000 4.425000 2.250000 ;
        RECT 4.350000 1.950000 4.725000 2.025000 ;
        RECT 4.425000 2.025000 4.650000 2.250000 ;
        RECT 4.425000 0.450000 4.650000 1.950000 ;
        RECT 4.650000 2.025000 4.725000 2.250000 ;
        RECT 7.650000 0.450000 7.950000 4.425000 ;
        RECT 7.575000 4.800000 8.025000 4.875000 ;
        RECT 7.575000 4.500000 7.650000 4.800000 ;
        RECT 7.575000 4.425000 8.025000 4.500000 ;
        RECT 7.650000 4.500000 7.950000 4.800000 ;
        RECT 7.950000 4.500000 8.025000 4.800000 ;
        END
        ANTENNADIFFAREA 0.708750 ;
    END GND
    OBS
        LAYER li1 ;
        RECT 1.050000 7.275000 6.225000 7.500000 ;
        RECT 1.050000 3.825000 1.275000 7.275000 ;
        RECT 1.050000 3.600000 1.575000 3.825000 ;
        RECT 1.575000 3.600000 1.875000 3.900000 ;
        RECT 1.500000 3.525000 1.950000 3.600000 ;
        RECT 1.500000 3.900000 1.950000 3.975000 ;
        RECT 1.500000 3.825000 1.575000 3.900000 ;
        RECT 1.875000 3.600000 1.950000 3.900000 ;
        RECT 3.000000 3.750000 3.225000 3.825000 ;
        RECT 3.000000 3.525000 3.225000 3.750000 ;
        RECT 3.000000 3.450000 3.225000 3.525000 ;
        RECT 3.600000 1.125000 3.975000 1.200000 ;
        RECT 3.600000 0.900000 3.675000 1.125000 ;
        RECT 3.600000 0.825000 3.975000 0.900000 ;
        RECT 3.675000 2.325000 3.750000 2.550000 ;
        RECT 3.675000 0.900000 3.900000 1.125000 ;
        RECT 3.750000 2.550000 3.975000 2.625000 ;
        RECT 3.750000 2.325000 3.975000 2.550000 ;
        RECT 3.750000 1.200000 3.975000 2.325000 ;
        RECT 3.900000 0.900000 6.150000 1.125000 ;
        RECT 5.025000 2.325000 5.325000 2.400000 ;
        RECT 5.025000 2.100000 5.100000 2.325000 ;
        RECT 5.025000 2.025000 5.400000 2.100000 ;
        RECT 5.100000 2.100000 5.325000 2.325000 ;
        RECT 5.325000 2.100000 5.400000 2.325000 ;
        RECT 5.850000 3.600000 6.225000 3.675000 ;
        RECT 5.850000 3.375000 5.925000 3.600000 ;
        RECT 5.850000 3.300000 6.225000 3.375000 ;
        RECT 6.000000 4.800000 6.225000 7.275000 ;
        RECT 5.925000 4.575000 6.225000 4.800000 ;
        RECT 5.925000 3.675000 6.150000 4.575000 ;
        RECT 5.925000 3.375000 6.150000 3.600000 ;
        RECT 6.150000 3.375000 6.225000 3.600000 ;
        RECT 6.075000 1.125000 6.525000 1.200000 ;
        RECT 6.600000 2.475000 6.975000 2.550000 ;
        RECT 6.075000 0.825000 6.150000 0.900000 ;
        RECT 6.075000 0.750000 6.525000 0.825000 ;
        RECT 6.150000 0.825000 6.450000 1.125000 ;
        RECT 6.450000 0.825000 6.525000 1.125000 ;
        RECT 6.600000 2.250000 6.675000 2.475000 ;
        RECT 6.600000 2.175000 6.975000 2.250000 ;
        RECT 6.675000 2.250000 6.900000 2.475000 ;
        RECT 6.900000 2.250000 6.975000 2.475000 ;
        LAYER met1 ;
        RECT 2.925000 3.750000 3.300000 3.825000 ;
        RECT 2.925000 3.525000 3.000000 3.750000 ;
        RECT 2.925000 3.450000 3.300000 3.525000 ;
        RECT 3.075000 1.200000 3.300000 3.450000 ;
        RECT 3.075000 1.125000 3.975000 1.200000 ;
        RECT 3.075000 0.900000 3.675000 1.125000 ;
        RECT 3.000000 3.525000 3.225000 3.750000 ;
        RECT 3.675000 0.900000 3.900000 1.125000 ;
        RECT 3.225000 3.525000 3.300000 3.750000 ;
        RECT 3.900000 0.900000 3.975000 1.125000 ;
        RECT 3.600000 0.825000 3.975000 0.900000 ;
        RECT 5.025000 2.325000 5.400000 2.400000 ;
        RECT 5.025000 2.100000 5.100000 2.325000 ;
        RECT 5.025000 2.025000 5.400000 2.100000 ;
        RECT 5.100000 2.100000 5.325000 2.325000 ;
        RECT 5.325000 2.250000 6.675000 2.325000 ;
        RECT 5.325000 2.175000 6.975000 2.250000 ;
        RECT 5.325000 2.100000 5.400000 2.175000 ;
        RECT 6.675000 2.250000 6.900000 2.475000 ;
        RECT 6.900000 2.250000 6.975000 2.475000 ;
        RECT 6.600000 2.475000 6.975000 2.550000 ;
        RECT 6.600000 2.325000 6.675000 2.475000 ;
    END
END _0_0std_0_0cells_0_0MUX2X1

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 2.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li1 ;
        RECT 0.600000 1.500000 0.900000 1.800000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li1 ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 445.800000 BY 448.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 445.800000 BY 448.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

