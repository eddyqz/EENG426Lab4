magic
tech sky130l
timestamp 1668303673
<< ndiffusion >>
rect 6 11 13 12
rect 6 8 7 11
rect 10 8 13 11
rect 6 6 13 8
rect 65 6 68 12
rect 70 11 77 12
rect 70 8 72 11
rect 75 8 77 11
rect 70 6 77 8
rect 79 6 82 12
rect 84 6 87 12
rect 89 10 94 12
rect 89 7 90 10
rect 93 7 94 10
rect 89 6 94 7
rect 98 11 105 12
rect 98 8 100 11
rect 103 8 105 11
rect 98 6 105 8
<< ndc >>
rect 7 8 10 11
rect 72 8 75 11
rect 90 7 93 10
rect 100 8 103 11
<< ntransistor >>
rect 13 6 65 12
rect 68 6 70 12
rect 77 6 79 12
rect 82 6 84 12
rect 87 6 89 12
rect 94 6 98 12
<< pdiffusion >>
rect 73 41 77 45
rect 8 39 13 41
rect 8 36 9 39
rect 12 36 13 39
rect 8 35 13 36
rect 51 35 68 41
rect 70 39 77 41
rect 70 36 72 39
rect 75 36 77 39
rect 70 35 77 36
rect 79 35 82 45
rect 84 35 87 45
rect 89 44 94 45
rect 89 41 90 44
rect 93 41 94 44
rect 89 35 94 41
rect 98 39 105 45
rect 98 36 100 39
rect 103 36 105 39
rect 98 35 105 36
<< pdc >>
rect 9 36 12 39
rect 72 36 75 39
rect 90 41 93 44
rect 100 36 103 39
<< ptransistor >>
rect 13 35 51 41
rect 68 35 70 41
rect 77 35 79 45
rect 82 35 84 45
rect 87 35 89 45
rect 94 35 98 45
<< polysilicon >>
rect 13 48 18 49
rect 13 45 14 48
rect 17 45 18 48
rect 77 45 79 47
rect 82 45 84 47
rect 87 45 89 47
rect 94 45 98 47
rect 13 43 18 45
rect 13 41 51 43
rect 68 41 70 43
rect 13 33 51 35
rect 68 26 70 35
rect 63 25 70 26
rect 63 22 64 25
rect 67 22 70 25
rect 63 21 70 22
rect 13 20 18 21
rect 13 17 14 20
rect 17 17 18 20
rect 13 14 18 17
rect 13 12 65 14
rect 68 12 70 21
rect 77 12 79 35
rect 82 12 84 35
rect 87 12 89 35
rect 94 26 98 35
rect 94 25 99 26
rect 94 22 95 25
rect 98 22 99 25
rect 94 21 99 22
rect 94 12 98 21
rect 13 4 65 6
rect 68 4 70 6
rect 77 -6 79 6
rect 72 -7 79 -6
rect 72 -11 73 -7
rect 77 -11 79 -7
rect 72 -12 79 -11
rect 82 -16 84 6
rect 87 -6 89 6
rect 94 4 98 6
rect 87 -7 97 -6
rect 87 -11 92 -7
rect 96 -11 97 -7
rect 87 -12 97 -11
rect 80 -17 86 -16
rect 80 -21 81 -17
rect 85 -21 86 -17
rect 80 -22 86 -21
<< pc >>
rect 14 45 17 48
rect 64 22 67 25
rect 14 17 17 20
rect 95 22 98 25
rect 73 -11 77 -7
rect 92 -11 96 -7
rect 81 -21 85 -17
<< m1 >>
rect 63 57 111 60
rect -9 48 18 49
rect -9 46 14 48
rect -9 22 -6 46
rect 13 45 14 46
rect 17 45 18 48
rect 13 44 18 45
rect 8 39 13 40
rect 8 36 9 39
rect 12 36 13 39
rect 8 35 13 36
rect 8 31 11 35
rect -1 30 11 31
rect -1 26 0 30
rect 4 28 11 30
rect 4 26 5 28
rect -1 25 5 26
rect -9 19 -3 22
rect -6 13 -3 19
rect 8 21 11 28
rect 63 26 66 57
rect 89 52 94 53
rect 89 49 90 52
rect 93 49 94 52
rect 89 48 94 49
rect 90 45 93 48
rect 89 44 94 45
rect 89 41 90 44
rect 93 41 94 44
rect 89 40 94 41
rect 71 39 76 40
rect 71 36 72 39
rect 75 36 76 39
rect 71 35 76 36
rect 99 39 104 40
rect 99 36 100 39
rect 103 36 104 39
rect 99 35 104 36
rect 108 35 111 57
rect 72 26 75 35
rect 99 33 111 35
rect 99 32 113 33
rect 99 31 108 32
rect 105 28 108 31
rect 112 28 113 32
rect 105 27 113 28
rect 63 25 68 26
rect 63 22 64 25
rect 67 22 68 25
rect 63 21 68 22
rect 72 25 99 26
rect 72 22 95 25
rect 98 22 99 25
rect 72 21 99 22
rect 8 20 18 21
rect 8 18 14 20
rect 13 17 14 18
rect 17 17 18 20
rect 13 16 18 17
rect -6 12 -1 13
rect 72 12 75 21
rect 105 16 108 27
rect 99 13 108 16
rect -6 9 -5 12
rect -2 11 11 12
rect -2 9 7 11
rect -6 8 7 9
rect 10 8 11 11
rect -6 0 -3 8
rect 6 7 11 8
rect 71 11 76 12
rect 99 11 104 13
rect 71 8 72 11
rect 75 8 76 11
rect 71 7 76 8
rect 89 10 94 11
rect 89 7 90 10
rect 93 7 94 10
rect 99 8 100 11
rect 103 8 104 11
rect 99 7 104 8
rect 89 6 94 7
rect 90 0 93 6
rect -6 -3 93 0
rect 72 -7 78 -6
rect 72 -11 73 -7
rect 77 -11 78 -7
rect 72 -12 78 -11
rect 91 -7 97 -6
rect 91 -11 92 -7
rect 96 -11 97 -7
rect 91 -12 97 -11
rect 80 -17 86 -16
rect 80 -21 81 -17
rect 85 -21 86 -17
rect 80 -22 86 -21
<< m2c >>
rect 0 26 4 30
rect 90 49 93 52
rect 108 28 112 32
rect -5 9 -2 12
<< m2 >>
rect -1 52 94 53
rect -1 50 90 52
rect -1 31 2 50
rect 89 49 90 50
rect 93 49 94 52
rect 89 48 94 49
rect 107 32 116 33
rect -1 30 5 31
rect -1 26 0 30
rect 4 26 5 30
rect 107 28 108 32
rect 112 28 116 32
rect 107 27 116 28
rect -1 25 5 26
rect -8 12 -1 13
rect -8 9 -5 12
rect -2 9 -1 12
rect -8 8 -1 9
<< labels >>
rlabel ndiffusion 99 7 99 7 3 #10
rlabel polysilicon 95 13 95 13 3 out
rlabel ndiffusion 90 7 90 7 3 GND
rlabel polysilicon 88 13 88 13 3 in(0)
rlabel polysilicon 83 13 83 13 3 in(1)
rlabel polysilicon 78 13 78 13 3 in(2)
rlabel ndiffusion 71 7 71 7 3 out
rlabel polysilicon 69 13 69 13 3 #10
rlabel polysilicon 14 13 14 13 3 Vdd
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 99 36 99 36 3 #10
rlabel polysilicon 95 34 95 34 3 out
rlabel pdiffusion 90 36 90 36 3 Vdd
rlabel polysilicon 88 34 88 34 3 in(0)
rlabel polysilicon 83 34 83 34 3 in(1)
rlabel polysilicon 78 34 78 34 3 in(2)
rlabel pdiffusion 71 36 71 36 3 out
rlabel polysilicon 69 34 69 34 3 #10
rlabel polysilicon 14 34 14 34 3 GND
rlabel pdiffusion 9 36 9 36 3 Vdd
rlabel m1 s 0 26 4 30 6 Vdd
port 5 nsew power input
rlabel m2c 1 27 1 27 3 Vdd
port 5 e
rlabel m1 0 9 0 9 3 GND
port 6 e
rlabel m1 s -1 8 3 12 6 GND
port 6 nsew ground input
rlabel m2c 109 29 109 29 3 out
port 4 e
rlabel m1 s 108 28 112 32 6 out
port 4 nsew signal output
rlabel m2 115 29 115 29 7 out
rlabel m2 -7 10 -7 10 3 GND
rlabel pc 93 -10 93 -10 3 in(0)
port 9 e
rlabel m1 s 92 -11 96 -7 6 in_50_6
port 1 nsew signal input
rlabel m1 s 81 -21 85 -17 6 in_51_6
port 2 nsew signal input
rlabel pc 82 -20 82 -20 3 in(1)
port 8 e
rlabel pc 74 -10 74 -10 3 in(2)
port 7 e
rlabel m1 s 73 -11 77 -7 6 in_52_6
port 3 nsew signal input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 112 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
