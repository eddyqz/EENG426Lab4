magic
tech sky130l
timestamp 1668326469
<< ndiffusion >>
rect 3 10 8 16
rect 3 7 4 10
rect 7 7 8 10
rect 3 6 8 7
rect 10 6 15 16
rect 17 10 22 16
rect 34 15 39 16
rect 34 12 35 15
rect 38 12 39 15
rect 34 10 39 12
rect 41 14 48 16
rect 41 11 43 14
rect 46 11 48 14
rect 41 10 48 11
rect 17 7 18 10
rect 21 7 22 10
rect 17 6 22 7
rect 44 6 48 10
rect 50 10 55 16
rect 50 7 51 10
rect 54 7 55 10
rect 50 6 55 7
rect 67 15 72 16
rect 67 12 68 15
rect 71 12 72 15
rect 67 6 72 12
rect 74 10 79 16
rect 74 7 75 10
rect 78 7 79 10
rect 74 6 79 7
<< ndc >>
rect 4 7 7 10
rect 35 12 38 15
rect 43 11 46 14
rect 18 7 21 10
rect 51 7 54 10
rect 68 12 71 15
rect 75 7 78 10
<< ntransistor >>
rect 8 6 10 16
rect 15 6 17 16
rect 39 10 41 16
rect 48 6 50 16
rect 72 6 74 16
<< pdiffusion >>
rect 3 47 8 48
rect 3 44 4 47
rect 7 44 8 47
rect 3 33 8 44
rect 10 41 14 48
rect 10 39 15 41
rect 10 36 11 39
rect 14 36 15 39
rect 10 33 15 36
rect 17 37 22 41
rect 17 34 18 37
rect 21 34 22 37
rect 17 33 22 34
rect 34 37 39 48
rect 34 34 35 37
rect 38 34 39 37
rect 34 33 39 34
rect 41 33 48 48
rect 50 37 55 48
rect 50 34 51 37
rect 54 34 55 37
rect 50 33 55 34
rect 67 47 72 48
rect 67 44 68 47
rect 71 44 72 47
rect 67 33 72 44
rect 74 37 79 48
rect 74 34 75 37
rect 78 34 79 37
rect 74 33 79 34
<< pdc >>
rect 4 44 7 47
rect 11 36 14 39
rect 18 34 21 37
rect 35 34 38 37
rect 51 34 54 37
rect 68 44 71 47
rect 75 34 78 37
<< ptransistor >>
rect 8 33 10 48
rect 15 33 17 41
rect 39 33 41 48
rect 48 33 50 48
rect 72 33 74 48
<< polysilicon >>
rect 72 57 77 58
rect 46 55 51 56
rect 15 52 23 53
rect 8 48 10 50
rect 15 49 19 52
rect 22 49 23 52
rect 15 48 23 49
rect 26 52 41 53
rect 26 49 27 52
rect 30 51 41 52
rect 46 52 47 55
rect 50 52 51 55
rect 46 51 51 52
rect 72 54 73 57
rect 76 54 77 57
rect 72 53 77 54
rect 30 49 31 51
rect 26 48 31 49
rect 39 48 41 51
rect 48 48 50 51
rect 72 48 74 53
rect 15 41 17 48
rect -1 25 4 26
rect 8 25 10 33
rect -1 22 0 25
rect 3 23 10 25
rect 3 22 4 23
rect -1 21 4 22
rect 8 16 10 23
rect 15 16 17 33
rect 39 16 41 33
rect 48 16 50 33
rect 72 16 74 33
rect 39 8 41 10
rect 8 4 10 6
rect 15 4 17 6
rect 48 4 50 6
rect 72 4 74 6
<< pc >>
rect 19 49 22 52
rect 27 49 30 52
rect 47 52 50 55
rect 73 54 76 57
rect 0 22 3 25
<< m1 >>
rect 63 68 68 69
rect 4 67 9 68
rect 4 64 5 67
rect 8 64 9 67
rect 63 65 64 68
rect 67 65 68 68
rect 63 64 68 65
rect 4 63 9 64
rect 4 47 7 63
rect 10 59 15 60
rect 10 56 11 59
rect 14 56 15 59
rect 10 55 15 56
rect 46 55 51 56
rect 4 43 7 44
rect 11 39 14 55
rect 18 52 23 53
rect 26 52 31 53
rect 18 49 19 52
rect 22 49 27 52
rect 30 49 31 52
rect 46 52 47 55
rect 50 52 51 55
rect 46 51 51 52
rect 18 48 23 49
rect 26 48 31 49
rect 64 48 67 64
rect 72 57 77 58
rect 72 54 73 57
rect 76 54 77 57
rect 72 53 77 54
rect 64 47 72 48
rect 64 44 68 47
rect 71 44 72 47
rect 67 43 72 44
rect 11 35 14 36
rect 18 37 21 38
rect 34 37 39 38
rect 18 33 21 34
rect 25 34 35 37
rect 38 34 39 37
rect 17 32 22 33
rect 17 29 18 32
rect 21 29 22 32
rect 17 28 22 29
rect -1 25 4 26
rect -1 22 0 25
rect 3 22 4 25
rect -1 21 4 22
rect 4 10 7 11
rect 4 3 7 7
rect 18 10 21 11
rect 25 10 28 34
rect 34 33 39 34
rect 50 37 60 38
rect 50 34 51 37
rect 54 34 56 37
rect 59 34 60 37
rect 50 33 60 34
rect 75 37 78 38
rect 78 34 85 37
rect 75 33 78 34
rect 33 20 38 21
rect 33 17 34 20
rect 37 17 38 20
rect 33 16 38 17
rect 35 15 38 16
rect 35 11 38 12
rect 43 14 46 15
rect 62 14 68 15
rect 62 11 63 14
rect 66 12 68 14
rect 71 12 72 15
rect 66 11 67 12
rect 21 7 28 10
rect 3 2 8 3
rect 3 -1 4 2
rect 7 -1 8 2
rect 3 -2 8 -1
rect 18 -6 21 7
rect 43 3 46 11
rect 51 10 54 11
rect 62 10 67 11
rect 75 10 78 11
rect 42 2 47 3
rect 42 -1 43 2
rect 46 -1 47 2
rect 51 2 54 7
rect 75 2 78 7
rect 51 -1 78 2
rect 42 -2 47 -1
rect 62 -6 67 -5
rect 82 -6 85 34
rect 18 -9 63 -6
rect 66 -9 85 -6
rect 18 -10 21 -9
rect 62 -10 67 -9
<< m2c >>
rect 5 64 8 67
rect 64 65 67 68
rect 11 56 14 59
rect 18 29 21 32
rect 56 34 59 37
rect 34 17 37 20
rect 63 11 66 14
rect 4 -1 7 2
rect 43 -1 46 2
rect 63 -9 66 -6
<< m2 >>
rect 63 68 68 69
rect 4 67 64 68
rect 4 64 5 67
rect 8 65 64 67
rect 67 65 68 68
rect 8 64 9 65
rect 63 64 68 65
rect 4 63 9 64
rect 10 59 15 60
rect 10 56 11 59
rect 14 56 59 59
rect 10 55 15 56
rect 56 38 59 56
rect 55 37 60 38
rect 55 34 56 37
rect 59 34 60 37
rect 55 33 60 34
rect 17 32 22 33
rect 17 29 18 32
rect 21 29 22 32
rect 17 28 22 29
rect 18 20 21 28
rect 33 20 38 21
rect 18 17 34 20
rect 37 17 38 20
rect 33 16 38 17
rect 62 14 67 15
rect 62 11 63 14
rect 66 11 67 14
rect 62 10 67 11
rect 3 2 8 3
rect 42 2 47 3
rect 3 -1 4 2
rect 7 -1 43 2
rect 46 -1 47 2
rect 3 -2 8 -1
rect 42 -2 47 -1
rect 63 -5 66 10
rect 62 -6 67 -5
rect 62 -9 63 -6
rect 66 -9 67 -6
rect 62 -10 67 -9
<< labels >>
rlabel ndiffusion 51 7 51 7 3 #10
rlabel polysilicon 49 17 49 17 3 B
rlabel ndiffusion 42 11 42 11 3 GND
rlabel polysilicon 40 17 40 17 3 S
rlabel ndiffusion 35 11 35 11 3 _S
rlabel polysilicon 49 32 49 32 3 B
rlabel pdiffusion 51 34 51 34 3 Vdd
rlabel polysilicon 40 32 40 32 3 S
rlabel pdiffusion 35 34 35 34 3 Y
rlabel ndiffusion 18 7 18 7 3 Y
rlabel polysilicon 16 17 16 17 3 S
rlabel polysilicon 9 17 9 17 3 A
rlabel ndiffusion 4 7 4 7 3 GND
rlabel pdiffusion 18 34 18 34 3 _S
rlabel polysilicon 16 32 16 32 3 S
rlabel pdiffusion 11 34 11 34 3 Vdd
rlabel polysilicon 9 32 9 32 3 A
rlabel pdiffusion 4 34 4 34 3 #5
rlabel ndiffusion 75 7 75 7 3 #10
rlabel polysilicon 73 17 73 17 3 _S
rlabel ndiffusion 68 7 68 7 3 Y
rlabel pdiffusion 75 34 75 34 3 Y
rlabel polysilicon 73 32 73 32 3 _S
rlabel pdiffusion 68 34 68 34 3 #5
rlabel m2 30 1 30 1 1 GND
rlabel m1 50 -8 50 -8 1 Y
rlabel m2 37 58 37 58 1 Vdd
rlabel m2 35 66 35 66 5 #5
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 80 48
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
