magic
tech sky130l
timestamp 1668317425
<< ndiffusion >>
rect 8 8 13 14
rect 8 5 9 8
rect 12 5 13 8
rect 8 4 13 5
rect 15 8 22 14
rect 15 5 17 8
rect 20 5 22 8
rect 15 4 22 5
rect 24 4 29 14
rect 25 -4 29 4
rect 31 8 36 14
rect 31 5 32 8
rect 35 5 36 8
rect 31 -4 36 5
rect 38 0 43 14
rect 38 -3 39 0
rect 42 -3 43 0
rect 38 -4 43 -3
rect 45 8 52 14
rect 45 5 46 8
rect 49 5 52 8
rect 45 -4 52 5
rect 48 -6 52 -4
rect 54 -2 59 14
rect 54 -5 55 -2
rect 58 -5 59 -2
rect 54 -6 59 -5
rect 61 -2 68 14
rect 61 -5 63 -2
rect 66 -5 68 -2
rect 61 -6 68 -5
rect 70 -2 75 14
rect 70 -5 71 -2
rect 74 -5 75 -2
rect 70 -6 75 -5
rect 77 13 84 14
rect 77 10 79 13
rect 82 10 84 13
rect 77 -6 84 10
rect 86 -6 89 14
rect 91 -6 94 14
rect 96 13 101 14
rect 96 10 97 13
rect 100 10 101 13
rect 96 8 101 10
rect 103 13 110 14
rect 103 10 106 13
rect 109 10 110 13
rect 103 8 110 10
rect 117 13 124 14
rect 117 10 118 13
rect 121 10 124 13
rect 117 8 124 10
rect 126 13 131 14
rect 126 10 127 13
rect 130 10 131 13
rect 126 8 131 10
rect 96 -6 100 8
<< ndc >>
rect 9 5 12 8
rect 17 5 20 8
rect 32 5 35 8
rect 39 -3 42 0
rect 46 5 49 8
rect 55 -5 58 -2
rect 63 -5 66 -2
rect 71 -5 74 -2
rect 79 10 82 13
rect 97 10 100 13
rect 106 10 109 13
rect 118 10 121 13
rect 127 10 130 13
<< ntransistor >>
rect 13 4 15 14
rect 22 4 24 14
rect 29 -4 31 14
rect 36 -4 38 14
rect 43 -4 45 14
rect 52 -6 54 14
rect 59 -6 61 14
rect 68 -6 70 14
rect 75 -6 77 14
rect 84 -6 86 14
rect 89 -6 91 14
rect 94 -6 96 14
rect 101 8 103 14
rect 124 8 126 14
<< pdiffusion >>
rect 64 67 68 71
rect 48 54 52 67
rect 18 42 22 54
rect 8 41 13 42
rect 8 38 9 41
rect 12 38 13 41
rect 8 31 13 38
rect 15 41 22 42
rect 15 38 17 41
rect 20 38 22 41
rect 15 31 22 38
rect 24 53 29 54
rect 24 50 25 53
rect 28 50 29 53
rect 24 31 29 50
rect 31 45 36 54
rect 31 42 32 45
rect 35 42 36 45
rect 31 31 36 42
rect 38 31 43 54
rect 45 53 52 54
rect 45 50 46 53
rect 49 50 52 53
rect 45 31 52 50
rect 54 66 59 67
rect 54 63 55 66
rect 58 63 59 66
rect 54 31 59 63
rect 61 61 68 67
rect 61 58 63 61
rect 66 58 68 61
rect 61 31 68 58
rect 70 67 74 71
rect 80 67 84 79
rect 70 66 75 67
rect 70 63 71 66
rect 74 63 75 66
rect 70 31 75 63
rect 77 35 84 67
rect 77 32 79 35
rect 82 32 84 35
rect 77 31 84 32
rect 86 31 89 79
rect 91 31 94 79
rect 96 39 100 79
rect 96 35 101 39
rect 96 32 97 35
rect 100 32 101 35
rect 96 31 101 32
rect 103 35 110 39
rect 103 32 106 35
rect 109 32 110 35
rect 103 31 110 32
rect 117 35 124 39
rect 117 32 118 35
rect 121 32 124 35
rect 117 31 124 32
rect 126 35 131 39
rect 126 32 127 35
rect 130 32 131 35
rect 126 31 131 32
<< pdc >>
rect 9 38 12 41
rect 17 38 20 41
rect 25 50 28 53
rect 32 42 35 45
rect 46 50 49 53
rect 55 63 58 66
rect 63 58 66 61
rect 71 63 74 66
rect 79 32 82 35
rect 97 32 100 35
rect 106 32 109 35
rect 118 32 121 35
rect 127 32 130 35
<< ptransistor >>
rect 13 31 15 42
rect 22 31 24 54
rect 29 31 31 54
rect 36 31 38 54
rect 43 31 45 54
rect 52 31 54 67
rect 59 31 61 67
rect 68 31 70 71
rect 75 31 77 67
rect 84 31 86 79
rect 89 31 91 79
rect 94 31 96 79
rect 101 31 103 39
rect 124 31 126 39
<< polysilicon >>
rect 22 131 24 136
rect 36 131 38 136
rect 52 131 54 136
rect 22 130 29 131
rect 22 127 25 130
rect 28 127 29 130
rect 22 126 29 127
rect 36 130 43 131
rect 36 127 39 130
rect 42 127 43 130
rect 36 126 43 127
rect 52 130 59 131
rect 52 127 55 130
rect 58 127 59 130
rect 52 126 59 127
rect 84 130 91 131
rect 84 127 85 130
rect 88 127 91 130
rect 84 126 91 127
rect 11 113 16 114
rect 11 110 12 113
rect 15 110 16 113
rect 11 109 16 110
rect 13 42 15 109
rect 22 54 24 126
rect 29 54 31 56
rect 36 54 38 126
rect 52 67 54 126
rect 59 114 61 119
rect 59 113 66 114
rect 59 110 62 113
rect 65 110 66 113
rect 59 109 66 110
rect 79 113 86 114
rect 79 110 80 113
rect 83 110 86 113
rect 79 109 86 110
rect 59 67 61 109
rect 84 79 86 109
rect 89 79 91 126
rect 94 79 96 81
rect 68 71 70 73
rect 43 54 45 56
rect 75 67 77 69
rect 101 39 103 41
rect 124 39 126 41
rect 13 29 15 31
rect 13 14 15 16
rect 22 14 24 31
rect 29 14 31 31
rect 36 14 38 31
rect 43 14 45 31
rect 52 14 54 31
rect 59 14 61 31
rect 68 14 70 31
rect 75 14 77 31
rect 84 14 86 31
rect 89 14 91 31
rect 94 14 96 31
rect 101 14 103 31
rect 124 14 126 31
rect 13 2 15 4
rect 22 2 24 4
rect 29 -56 31 -4
rect 36 -6 38 -4
rect 43 -56 45 -4
rect 101 6 103 8
rect 124 6 126 8
rect 101 5 109 6
rect 101 2 105 5
rect 108 2 109 5
rect 101 1 109 2
rect 124 5 130 6
rect 124 2 126 5
rect 129 2 130 5
rect 124 1 130 2
rect 52 -8 54 -6
rect 59 -8 61 -6
rect 68 -18 70 -6
rect 75 -18 77 -6
rect 84 -8 86 -6
rect 89 -8 91 -6
rect 68 -19 77 -18
rect 68 -22 71 -19
rect 74 -22 77 -19
rect 68 -23 77 -22
rect 68 -56 70 -23
rect 94 -56 96 -6
rect 29 -57 36 -56
rect 29 -60 32 -57
rect 35 -60 36 -57
rect 29 -61 36 -60
rect 43 -57 50 -56
rect 43 -60 46 -57
rect 49 -60 50 -57
rect 43 -61 50 -60
rect 68 -57 75 -56
rect 68 -60 71 -57
rect 74 -60 75 -57
rect 68 -61 75 -60
rect 89 -57 96 -56
rect 89 -60 90 -57
rect 93 -60 96 -57
rect 89 -61 96 -60
<< pc >>
rect 25 127 28 130
rect 39 127 42 130
rect 55 127 58 130
rect 85 127 88 130
rect 12 110 15 113
rect 62 110 65 113
rect 80 110 83 113
rect 105 2 108 5
rect 126 2 129 5
rect 71 -22 74 -19
rect 32 -60 35 -57
rect 46 -60 49 -57
rect 71 -60 74 -57
rect 90 -60 93 -57
<< m1 >>
rect 24 135 29 136
rect 24 132 25 135
rect 28 132 29 135
rect 24 130 29 132
rect 24 127 25 130
rect 28 127 29 130
rect 24 126 29 127
rect 38 135 43 136
rect 38 132 39 135
rect 42 132 43 135
rect 38 130 43 132
rect 38 127 39 130
rect 42 127 43 130
rect 38 126 43 127
rect 54 135 59 136
rect 54 132 55 135
rect 58 132 59 135
rect 54 130 59 132
rect 54 127 55 130
rect 58 127 59 130
rect 54 126 59 127
rect 84 135 89 136
rect 84 132 85 135
rect 88 132 89 135
rect 84 130 89 132
rect 84 127 85 130
rect 88 127 89 130
rect 84 126 89 127
rect 11 118 16 119
rect 11 115 12 118
rect 15 115 16 118
rect 11 113 16 115
rect 11 110 12 113
rect 15 110 16 113
rect 11 109 16 110
rect 61 118 66 119
rect 61 115 62 118
rect 65 115 66 118
rect 61 113 66 115
rect 61 110 62 113
rect 65 110 66 113
rect 61 109 66 110
rect 79 118 84 119
rect 79 115 80 118
rect 83 115 84 118
rect 79 113 84 115
rect 79 110 80 113
rect 83 110 84 113
rect 79 109 84 110
rect 45 100 50 101
rect 45 97 46 100
rect 49 97 50 100
rect 45 96 50 97
rect 96 100 101 101
rect 96 97 97 100
rect 100 97 101 100
rect 96 96 101 97
rect 46 82 49 96
rect 54 90 59 91
rect 54 87 55 90
rect 58 87 59 90
rect 54 86 59 87
rect 70 90 75 91
rect 70 87 71 90
rect 74 87 75 90
rect 70 86 75 87
rect 8 81 13 82
rect 8 78 9 81
rect 12 78 13 81
rect 8 77 13 78
rect 45 81 50 82
rect 45 78 46 81
rect 49 78 50 81
rect 45 77 50 78
rect 9 42 12 77
rect 24 72 29 73
rect 24 69 25 72
rect 28 69 29 72
rect 24 68 29 69
rect 16 62 21 63
rect 16 59 17 62
rect 20 59 21 62
rect 16 58 21 59
rect 17 42 20 58
rect 25 54 28 68
rect 31 62 36 63
rect 31 59 32 62
rect 35 59 36 62
rect 31 58 36 59
rect 24 53 29 54
rect 24 50 25 53
rect 28 50 29 53
rect 24 49 29 50
rect 32 46 35 58
rect 46 54 49 77
rect 55 67 58 86
rect 62 81 67 82
rect 62 78 63 81
rect 66 78 67 81
rect 62 77 67 78
rect 54 66 59 67
rect 54 63 55 66
rect 58 63 59 66
rect 54 62 59 63
rect 63 62 66 77
rect 71 67 74 86
rect 70 66 75 67
rect 70 63 71 66
rect 74 63 75 66
rect 70 62 75 63
rect 62 61 67 62
rect 62 58 63 61
rect 66 58 67 61
rect 62 57 67 58
rect 45 53 50 54
rect 45 50 46 53
rect 49 50 50 53
rect 45 49 50 50
rect 97 50 100 96
rect 117 57 122 58
rect 135 57 140 58
rect 117 54 118 57
rect 121 54 136 57
rect 139 54 140 57
rect 117 53 122 54
rect 135 53 140 54
rect 97 49 105 50
rect 97 46 101 49
rect 104 46 105 49
rect 31 45 36 46
rect 31 42 32 45
rect 35 42 36 45
rect 8 41 13 42
rect 8 38 9 41
rect 12 38 13 41
rect 8 37 13 38
rect 16 41 21 42
rect 31 41 36 42
rect 97 45 105 46
rect 16 38 17 41
rect 20 38 21 41
rect 16 37 21 38
rect 97 36 100 45
rect 118 36 121 53
rect 126 49 131 50
rect 126 46 127 49
rect 130 46 131 49
rect 126 45 131 46
rect 127 36 130 45
rect 78 35 83 36
rect 78 32 79 35
rect 82 32 83 35
rect 78 31 83 32
rect 96 35 101 36
rect 96 32 97 35
rect 100 32 101 35
rect 96 31 101 32
rect 105 35 110 36
rect 105 32 106 35
rect 109 32 110 35
rect 105 31 110 32
rect 117 35 122 36
rect 117 32 118 35
rect 121 32 122 35
rect 117 31 122 32
rect 126 35 131 36
rect 126 32 127 35
rect 130 32 131 35
rect 126 31 131 32
rect 79 14 82 31
rect 106 14 109 31
rect 78 13 83 14
rect 78 10 79 13
rect 82 10 83 13
rect 78 9 83 10
rect 96 13 101 14
rect 96 10 97 13
rect 100 10 101 13
rect 96 9 101 10
rect 105 13 110 14
rect 105 10 106 13
rect 109 10 110 13
rect 105 9 110 10
rect 117 13 122 14
rect 117 10 118 13
rect 121 10 122 13
rect 117 9 122 10
rect 126 13 131 14
rect 136 13 139 53
rect 126 10 127 13
rect 130 10 139 13
rect 126 9 131 10
rect 8 8 13 9
rect 8 5 9 8
rect 12 5 13 8
rect 8 4 13 5
rect 16 8 21 9
rect 16 5 17 8
rect 20 5 21 8
rect 16 4 21 5
rect 31 8 36 9
rect 31 5 32 8
rect 35 5 36 8
rect 31 4 36 5
rect 45 8 50 9
rect 45 5 46 8
rect 49 5 50 8
rect 45 4 50 5
rect 9 -10 12 4
rect 17 1 20 4
rect 16 0 21 1
rect 16 -3 17 0
rect 20 -3 21 0
rect 16 -4 21 -3
rect 8 -11 13 -10
rect 8 -14 9 -11
rect 12 -14 13 -11
rect 8 -15 13 -14
rect 17 -42 20 -4
rect 32 -19 35 4
rect 38 0 43 1
rect 38 -3 39 0
rect 42 -3 43 0
rect 38 -4 43 -3
rect 39 -10 42 -4
rect 38 -11 43 -10
rect 38 -14 39 -11
rect 42 -14 43 -11
rect 38 -15 43 -14
rect 46 -19 49 4
rect 54 -2 59 -1
rect 54 -5 55 -2
rect 58 -5 59 -2
rect 54 -6 59 -5
rect 62 -2 67 -1
rect 62 -5 63 -2
rect 66 -5 67 -2
rect 62 -6 67 -5
rect 70 -2 75 -1
rect 70 -5 71 -2
rect 74 -5 75 -2
rect 70 -6 75 -5
rect 55 -10 58 -6
rect 54 -11 59 -10
rect 54 -14 55 -11
rect 58 -14 59 -11
rect 54 -15 59 -14
rect 31 -20 36 -19
rect 31 -23 32 -20
rect 35 -23 36 -20
rect 31 -24 36 -23
rect 45 -20 50 -19
rect 45 -23 46 -20
rect 49 -23 50 -20
rect 45 -24 50 -23
rect 46 -29 49 -24
rect 63 -29 66 -6
rect 71 -10 74 -6
rect 70 -11 75 -10
rect 70 -14 71 -11
rect 74 -14 75 -11
rect 70 -15 75 -14
rect 70 -19 75 -18
rect 70 -22 71 -19
rect 74 -22 75 -19
rect 70 -24 75 -22
rect 79 -24 82 9
rect 97 -14 100 9
rect 104 5 109 6
rect 104 2 105 5
rect 108 2 109 5
rect 104 1 109 2
rect 96 -15 101 -14
rect 96 -18 97 -15
rect 100 -18 101 -15
rect 96 -19 101 -18
rect 70 -27 71 -24
rect 74 -27 75 -24
rect 70 -28 75 -27
rect 78 -25 83 -24
rect 78 -28 79 -25
rect 82 -28 83 -25
rect 78 -29 83 -28
rect 45 -30 50 -29
rect 45 -33 46 -30
rect 49 -33 50 -30
rect 45 -34 50 -33
rect 62 -30 67 -29
rect 62 -33 63 -30
rect 66 -33 67 -30
rect 62 -34 67 -33
rect 46 -37 49 -34
rect 97 -37 100 -19
rect 105 -31 108 1
rect 118 -14 121 9
rect 125 5 130 6
rect 125 2 126 5
rect 129 2 130 5
rect 125 1 130 2
rect 117 -15 122 -14
rect 117 -18 118 -15
rect 121 -18 122 -15
rect 117 -19 122 -18
rect 126 -24 129 1
rect 125 -25 130 -24
rect 125 -28 126 -25
rect 129 -28 130 -25
rect 125 -29 130 -28
rect 104 -32 109 -31
rect 104 -35 105 -32
rect 108 -35 109 -32
rect 104 -36 109 -35
rect 45 -38 50 -37
rect 45 -41 46 -38
rect 49 -41 50 -38
rect 45 -42 50 -41
rect 96 -38 101 -37
rect 96 -41 97 -38
rect 100 -41 101 -38
rect 96 -42 101 -41
rect 16 -43 21 -42
rect 16 -46 17 -43
rect 20 -46 21 -43
rect 16 -47 21 -46
rect 31 -52 36 -51
rect 31 -55 32 -52
rect 35 -55 36 -52
rect 31 -57 36 -55
rect 31 -60 32 -57
rect 35 -60 36 -57
rect 31 -61 36 -60
rect 45 -52 50 -51
rect 45 -55 46 -52
rect 49 -55 50 -52
rect 45 -57 50 -55
rect 45 -60 46 -57
rect 49 -60 50 -57
rect 45 -61 50 -60
rect 70 -52 75 -51
rect 70 -55 71 -52
rect 74 -55 75 -52
rect 70 -57 75 -55
rect 70 -60 71 -57
rect 74 -60 75 -57
rect 70 -61 75 -60
rect 89 -52 94 -51
rect 89 -55 90 -52
rect 93 -55 94 -52
rect 89 -57 94 -55
rect 89 -60 90 -57
rect 93 -60 94 -57
rect 89 -61 94 -60
<< m2c >>
rect 25 132 28 135
rect 39 132 42 135
rect 55 132 58 135
rect 85 132 88 135
rect 12 115 15 118
rect 62 115 65 118
rect 80 115 83 118
rect 46 97 49 100
rect 97 97 100 100
rect 55 87 58 90
rect 71 87 74 90
rect 9 78 12 81
rect 46 78 49 81
rect 25 69 28 72
rect 17 59 20 62
rect 32 59 35 62
rect 63 78 66 81
rect 118 54 121 57
rect 136 54 139 57
rect 101 46 104 49
rect 127 46 130 49
rect 17 -3 20 0
rect 9 -14 12 -11
rect 39 -14 42 -11
rect 55 -14 58 -11
rect 32 -23 35 -20
rect 46 -23 49 -20
rect 71 -14 74 -11
rect 97 -18 100 -15
rect 71 -27 74 -24
rect 79 -28 82 -25
rect 46 -33 49 -30
rect 63 -33 66 -30
rect 118 -18 121 -15
rect 126 -28 129 -25
rect 105 -35 108 -32
rect 46 -41 49 -38
rect 97 -41 100 -38
rect 17 -46 20 -43
rect 32 -55 35 -52
rect 46 -55 49 -52
rect 71 -55 74 -52
rect 90 -55 93 -52
<< m2 >>
rect 24 135 29 136
rect 38 135 43 136
rect 54 135 59 136
rect 84 135 89 136
rect 24 132 25 135
rect 28 132 39 135
rect 42 132 55 135
rect 58 132 85 135
rect 88 132 89 135
rect 24 131 29 132
rect 38 131 43 132
rect 54 131 59 132
rect 84 131 89 132
rect 11 118 16 119
rect 61 118 66 119
rect 79 118 84 119
rect 11 115 12 118
rect 15 115 62 118
rect 65 115 80 118
rect 83 115 84 118
rect 11 114 16 115
rect 61 114 66 115
rect 79 114 84 115
rect 45 100 50 101
rect 96 100 101 101
rect 45 97 46 100
rect 49 97 97 100
rect 100 97 101 100
rect 45 96 50 97
rect 96 96 101 97
rect 54 90 59 91
rect 70 90 75 91
rect 54 87 55 90
rect 58 87 71 90
rect 74 87 75 90
rect 54 86 59 87
rect 70 86 75 87
rect 8 81 13 82
rect 45 81 50 82
rect 62 81 67 82
rect 8 78 9 81
rect 12 78 46 81
rect 49 78 63 81
rect 66 78 67 81
rect 8 77 13 78
rect 45 77 50 78
rect 62 77 67 78
rect 24 72 29 73
rect 2 69 25 72
rect 28 69 29 72
rect 2 0 5 69
rect 24 68 29 69
rect 16 62 21 63
rect 31 62 36 63
rect 16 59 17 62
rect 20 59 32 62
rect 35 59 36 62
rect 16 58 21 59
rect 31 58 36 59
rect 117 57 122 58
rect 117 54 118 57
rect 121 54 122 57
rect 117 53 122 54
rect 135 57 140 58
rect 135 54 136 57
rect 139 54 140 57
rect 135 53 140 54
rect 100 49 105 50
rect 126 49 131 50
rect 100 46 101 49
rect 104 46 127 49
rect 130 46 131 49
rect 100 45 105 46
rect 126 45 131 46
rect 16 0 21 1
rect 2 -3 17 0
rect 20 -3 21 0
rect 16 -4 21 -3
rect 8 -11 13 -10
rect 38 -11 43 -10
rect 8 -14 9 -11
rect 12 -14 39 -11
rect 42 -14 43 -11
rect 8 -15 13 -14
rect 38 -15 43 -14
rect 54 -11 59 -10
rect 70 -11 75 -10
rect 54 -14 55 -11
rect 58 -14 71 -11
rect 74 -14 75 -11
rect 54 -15 59 -14
rect 70 -15 75 -14
rect 96 -15 101 -14
rect 117 -15 122 -14
rect 96 -18 97 -15
rect 100 -18 118 -15
rect 121 -18 122 -15
rect 96 -19 101 -18
rect 117 -19 122 -18
rect 31 -20 36 -19
rect 45 -20 50 -19
rect 31 -23 32 -20
rect 35 -23 46 -20
rect 49 -23 50 -20
rect 31 -24 36 -23
rect 45 -24 50 -23
rect 70 -24 75 -23
rect 70 -27 71 -24
rect 74 -27 75 -24
rect 70 -28 75 -27
rect 78 -25 83 -24
rect 125 -25 130 -24
rect 78 -28 79 -25
rect 82 -28 126 -25
rect 129 -28 130 -25
rect 45 -30 50 -29
rect 62 -30 67 -29
rect 45 -33 46 -30
rect 49 -33 63 -30
rect 66 -33 67 -30
rect 45 -34 50 -33
rect 62 -34 67 -33
rect 71 -31 74 -28
rect 78 -29 83 -28
rect 125 -29 130 -28
rect 71 -32 109 -31
rect 71 -34 105 -32
rect 104 -35 105 -34
rect 108 -35 109 -32
rect 104 -36 109 -35
rect 45 -38 50 -37
rect 96 -38 101 -37
rect 45 -41 46 -38
rect 49 -41 97 -38
rect 100 -41 101 -38
rect 45 -42 50 -41
rect 96 -42 101 -41
rect 16 -43 21 -42
rect 16 -46 17 -43
rect 20 -44 21 -43
rect 105 -44 108 -36
rect 20 -46 108 -44
rect 16 -47 108 -46
rect 31 -52 36 -51
rect 31 -55 32 -52
rect 35 -55 36 -52
rect 31 -56 36 -55
rect 45 -52 50 -51
rect 45 -55 46 -52
rect 49 -55 50 -52
rect 45 -56 50 -55
rect 70 -52 75 -51
rect 70 -55 71 -52
rect 74 -55 75 -52
rect 70 -56 75 -55
rect 89 -52 94 -51
rect 89 -55 90 -52
rect 93 -55 94 -52
rect 89 -56 94 -55
<< labels >>
rlabel pdiffusion 104 32 104 32 3 YC
rlabel pdiffusion 97 32 97 32 3 Vdd
rlabel polysilicon 102 30 102 30 3 _YC
rlabel polysilicon 95 30 95 30 3 A
rlabel polysilicon 90 30 90 30 3 B
rlabel pdiffusion 78 32 78 32 3 _YS
rlabel polysilicon 85 30 85 30 3 C
rlabel pdiffusion 71 32 71 32 3 #12
rlabel polysilicon 76 30 76 30 3 _YC
rlabel polysilicon 69 30 69 30 3 A
rlabel pdiffusion 62 32 62 32 3 Vdd
rlabel polysilicon 60 30 60 30 3 C
rlabel pdiffusion 55 32 55 32 3 #12
rlabel polysilicon 53 30 53 30 3 B
rlabel pdiffusion 46 32 46 32 3 Vdd
rlabel polysilicon 44 30 44 30 3 A
rlabel polysilicon 37 30 37 30 3 B
rlabel pdiffusion 32 32 32 32 3 #8
rlabel polysilicon 30 30 30 30 3 A
rlabel pdiffusion 25 32 25 32 3 _YC
rlabel polysilicon 23 30 23 30 3 B
rlabel pdiffusion 16 32 16 32 3 #8
rlabel polysilicon 14 30 14 30 3 C
rlabel pdiffusion 9 32 9 32 3 Vdd
rlabel polysilicon 102 15 102 15 3 _YC
rlabel polysilicon 95 15 95 15 3 A
rlabel polysilicon 90 15 90 15 3 B
rlabel polysilicon 85 15 85 15 3 C
rlabel ndiffusion 104 9 104 9 3 YC
rlabel polysilicon 76 15 76 15 3 _YC
rlabel ndiffusion 97 -5 97 -5 3 GND
rlabel polysilicon 69 15 69 15 3 A
rlabel polysilicon 60 15 60 15 3 C
rlabel polysilicon 53 15 53 15 3 B
rlabel ndiffusion 78 -5 78 -5 3 _YS
rlabel ndiffusion 46 5 46 5 3 GND
rlabel polysilicon 44 15 44 15 3 A
rlabel ndiffusion 71 -5 71 -5 3 #15
rlabel polysilicon 37 15 37 15 3 B
rlabel ndiffusion 62 -5 62 -5 3 GND
rlabel ndiffusion 32 5 32 5 3 GND
rlabel polysilicon 30 15 30 15 3 A
rlabel ndiffusion 55 -5 55 -5 3 #15
rlabel polysilicon 23 15 23 15 3 B
rlabel ndiffusion 16 5 16 5 3 _YC
rlabel polysilicon 14 15 14 15 3 C
rlabel ndiffusion 9 5 9 5 3 #3
rlabel pdiffusion 127 32 127 32 3 Vdd
rlabel polysilicon 125 30 125 30 3 _YS
rlabel pdiffusion 120 32 120 32 3 YS
rlabel ndiffusion 127 9 127 9 3 YS
rlabel polysilicon 125 15 125 15 3 _YS
rlabel ndiffusion 120 9 120 9 3 GND
rlabel m2 26 -13 26 -13 1 #3
rlabel m2 39 -21 39 -21 1 GND
rlabel m2 70 -39 70 -39 1 GND
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 144 88
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
