magic
tech sky130l
timestamp 1668328199
<< error_p >>
rect 24 13 25 15
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 8 12 11
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 24 13 29
rect 8 21 9 24
rect 12 21 13 24
rect 8 19 13 21
rect 15 24 20 29
rect 15 21 16 24
rect 19 21 20 24
rect 15 19 20 21
<< pdc >>
rect 9 21 12 24
rect 16 21 19 24
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 29 15 31
rect 13 17 15 19
rect 24 17 29 18
rect 13 15 25 17
rect 13 12 15 15
rect 24 14 25 15
rect 28 14 29 17
rect 24 13 29 14
rect 13 4 15 6
<< pc >>
rect 25 14 28 17
<< m1 >>
rect 3 24 13 25
rect 3 21 4 24
rect 7 21 9 24
rect 12 21 13 24
rect 3 20 13 21
rect 16 24 19 25
rect 19 21 28 24
rect 16 20 19 21
rect 25 18 28 21
rect 24 17 29 18
rect 24 14 25 17
rect 28 14 29 17
rect 24 13 29 14
rect 3 11 13 12
rect 3 8 4 11
rect 7 8 9 11
rect 12 8 13 11
rect 3 7 13 8
rect 16 11 22 12
rect 19 8 22 11
rect 16 7 22 8
<< m2c >>
rect 4 21 7 24
rect 4 8 7 11
<< m2 >>
rect 1 24 8 25
rect 1 21 4 24
rect 7 21 8 24
rect 1 20 8 21
rect 1 11 8 12
rect 1 8 4 11
rect 7 8 8 11
rect 1 7 8 8
<< labels >>
rlabel ndiffusion 16 7 16 7 3 Y
rlabel pdiffusion 16 20 16 20 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel polysilicon 14 18 14 18 3 x
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m2 2 9 2 9 2 GND
rlabel m2 2 23 2 23 3 Vdd
rlabel m1 26 22 26 22 7 x
rlabel m1 21 9 21 9 1 Y
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 32 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
