magic
tech sky130l
timestamp 1668573647
<< ndiffusion >>
rect 16 14 21 16
rect 16 11 17 14
rect 20 11 21 14
rect 16 10 21 11
rect 23 14 28 16
rect 23 11 24 14
rect 27 11 28 14
rect 23 10 28 11
rect 30 14 35 16
rect 30 11 31 14
rect 34 11 35 14
rect 30 10 35 11
<< ndc >>
rect 17 11 20 14
rect 24 11 27 14
rect 31 11 34 14
<< ntransistor >>
rect 21 10 23 16
rect 28 10 30 16
<< pdiffusion >>
rect 16 32 21 38
rect 16 29 17 32
rect 20 29 21 32
rect 16 23 21 29
rect 23 23 28 38
rect 30 32 35 38
rect 30 29 31 32
rect 34 29 35 32
rect 30 23 35 29
<< pdc >>
rect 17 29 20 32
rect 31 29 34 32
<< ptransistor >>
rect 21 23 23 38
rect 28 23 30 38
<< polysilicon >>
rect 15 45 20 46
rect 15 42 16 45
rect 19 42 20 45
rect 15 41 20 42
rect 26 45 31 46
rect 26 42 27 45
rect 30 42 31 45
rect 26 41 31 42
rect 16 39 23 41
rect 21 38 23 39
rect 28 38 30 41
rect 21 16 23 23
rect 28 16 30 23
rect 21 8 23 10
rect 28 8 30 10
<< pc >>
rect 16 42 19 45
rect 27 42 30 45
<< m1 >>
rect 7 41 12 47
rect 15 45 20 47
rect 15 42 16 45
rect 19 42 20 45
rect 15 41 20 42
rect 26 45 31 47
rect 26 42 27 45
rect 30 42 31 45
rect 35 43 44 47
rect 26 41 31 42
rect 7 38 8 41
rect 11 38 12 41
rect 7 32 12 38
rect 31 32 34 33
rect 7 29 17 32
rect 20 29 21 32
rect 7 2 12 29
rect 31 21 34 29
rect 24 18 34 21
rect 16 14 21 15
rect 16 11 17 14
rect 20 11 21 14
rect 16 10 21 11
rect 24 14 27 18
rect 39 14 44 43
rect 30 11 31 14
rect 34 11 40 14
rect 43 11 44 14
rect 15 6 20 7
rect 15 3 16 6
rect 19 5 20 6
rect 24 5 27 11
rect 39 5 44 11
rect 19 3 27 5
rect 15 2 27 3
rect 31 2 44 5
<< m2c >>
rect 16 42 19 45
rect 27 42 30 45
rect 8 38 11 41
rect 17 11 20 14
rect 40 11 43 14
rect 16 3 19 6
<< m2 >>
rect 15 45 20 46
rect 15 42 16 45
rect 19 42 20 45
rect 7 41 12 42
rect 15 41 20 42
rect 26 45 31 46
rect 26 42 27 45
rect 30 42 31 45
rect 26 41 31 42
rect 7 38 8 41
rect 11 38 12 41
rect 7 37 12 38
rect 16 14 44 15
rect 16 11 17 14
rect 20 11 40 14
rect 43 11 44 14
rect 16 10 44 11
rect 15 6 20 7
rect 15 3 16 6
rect 19 3 20 6
rect 15 2 20 3
<< labels >>
rlabel polysilicon 29 39 29 39 3 B
rlabel ndiffusion 28 12 28 12 3 Y
rlabel pdiffusion 31 24 31 24 3 Y
rlabel polysilicon 29 9 29 9 3 B
rlabel ntransistor 29 11 29 11 3 B
rlabel polysilicon 29 17 29 17 3 B
rlabel ptransistor 29 24 29 24 3 B
rlabel polysilicon 22 39 22 39 3 A
rlabel polysilicon 22 17 22 17 3 A
rlabel ptransistor 22 24 22 24 3 A
rlabel pdiffusion 17 24 17 24 3 Vdd
rlabel polysilicon 17 40 17 40 3 A
rlabel m1 32 22 32 22 3 Y
port 1 e
rlabel ndc 25 12 25 12 3 Y
port 1 e
rlabel pc 28 43 28 43 3 B
port 2 e
rlabel m1 27 42 27 42 3 B
port 2 e
rlabel m1 27 43 27 43 3 B
port 2 e
rlabel m1 27 46 27 46 3 B
port 2 e
rlabel m1 25 6 25 6 3 Y
port 1 e
rlabel m1 25 15 25 15 3 Y
port 1 e
rlabel m1 25 19 25 19 3 Y
port 1 e
rlabel pc 17 43 17 43 3 A
port 3 e
rlabel m1 16 42 16 42 3 A
port 3 e
rlabel m1 16 43 16 43 3 A
port 3 e
rlabel m1 16 46 16 46 3 A
port 3 e
rlabel m1 17 3 17 3 3 Y
port 1 e
rlabel m1 15 30 15 30 1 Vdd
rlabel m2c 10 39 10 39 3 Vdd
rlabel m2c 42 13 42 13 7 GND
rlabel m2c 18 12 18 12 1 GND
rlabel pdc 33 30 33 30 1 Y
rlabel m1 42 32 42 32 7 GND
rlabel m1 8 26 8 26 3 Vdd
rlabel m1 10 6 10 6 2 Vdd
<< end >>
