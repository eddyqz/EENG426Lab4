magic
tech sky130l
timestamp 1668469005
<< checkpaint >>
rect -24 78 61 80
rect -24 72 62 78
rect -24 66 68 72
rect -26 -3 68 66
rect -24 -19 68 -3
rect -24 -22 59 -19
rect -19 -24 59 -22
rect -10 -28 59 -24
<< ndiffusion >>
rect 8 17 13 20
rect 8 14 9 17
rect 12 14 13 17
rect 8 10 13 14
rect 15 10 20 20
rect 22 10 27 20
<< ndc >>
rect 9 14 12 17
<< ntransistor >>
rect 13 10 15 20
rect 20 10 22 20
<< pdiffusion >>
rect 8 33 13 35
rect 8 30 9 33
rect 12 30 13 33
rect 8 27 13 30
rect 15 32 20 35
rect 15 29 16 32
rect 19 29 20 32
rect 15 27 20 29
rect 22 32 27 35
rect 22 29 23 32
rect 26 29 27 32
rect 22 27 27 29
<< pdc >>
rect 9 30 12 33
rect 16 29 19 32
rect 23 29 26 32
<< ptransistor >>
rect 13 27 15 35
rect 20 27 22 35
<< polysilicon >>
rect 8 46 13 47
rect 8 43 9 46
rect 12 43 13 46
rect 8 38 13 43
rect 18 46 23 47
rect 18 43 19 46
rect 22 43 23 46
rect 8 36 15 38
rect 18 36 23 43
rect 13 35 15 36
rect 20 35 22 36
rect 13 20 15 27
rect 20 20 22 27
rect 13 8 15 10
rect 20 8 22 10
<< pc >>
rect 9 43 12 46
rect 19 43 22 46
<< m1 >>
rect 8 46 13 48
rect 8 43 9 46
rect 12 43 13 46
rect 18 46 23 48
rect 18 43 19 46
rect 22 43 23 46
rect 26 45 29 48
rect 8 37 12 43
rect 18 36 22 43
rect 6 33 13 34
rect 6 30 9 33
rect 12 30 13 33
rect 6 29 13 30
rect 16 32 19 33
rect 22 29 23 32
rect 26 29 29 42
rect 16 25 19 29
rect 16 21 27 25
rect 8 17 13 18
rect 8 14 9 17
rect 12 14 13 17
rect 8 13 13 14
rect 22 4 27 21
rect 32 17 36 40
rect 35 14 36 17
rect 32 13 36 14
<< m2c >>
rect 26 42 29 45
rect 9 30 12 33
rect 9 14 12 17
rect 32 14 35 17
<< m2 >>
rect 25 45 30 46
rect 25 42 26 45
rect 29 42 30 45
rect 25 34 30 42
rect 8 33 30 34
rect 8 30 9 33
rect 12 30 30 33
rect 8 29 30 30
rect 8 17 36 18
rect 8 14 9 17
rect 12 14 32 17
rect 35 14 36 17
rect 8 13 36 14
<< labels >>
rlabel ndiffusion 23 11 23 11 3 Y
rlabel pdiffusion 23 28 23 28 3 Vdd
rlabel pdiffusion 23 33 23 33 3 Vdd
rlabel pdiffusion 20 30 20 30 3 Y
rlabel polysilicon 21 36 21 36 3 B
rlabel polysilicon 21 9 21 9 3 B
rlabel ntransistor 21 11 21 11 3 B
rlabel polysilicon 21 21 21 21 3 B
rlabel ptransistor 21 28 21 28 3 B
rlabel pdiffusion 16 28 16 28 3 Y
rlabel pdiffusion 16 30 16 30 3 Y
rlabel pdiffusion 16 33 16 33 3 Y
rlabel polysilicon 14 9 14 9 3 A
rlabel ntransistor 14 11 14 11 3 A
rlabel polysilicon 14 21 14 21 3 A
rlabel ptransistor 14 28 14 28 3 A
rlabel polysilicon 14 36 14 36 3 A
rlabel ndiffusion 9 11 9 11 3 GND
rlabel pdiffusion 9 28 9 28 3 Vdd
rlabel polysilicon 9 37 9 37 3 A
rlabel polysilicon 9 39 9 39 3 A
rlabel m1 27 30 27 30 3 Vdd
rlabel m1 27 46 27 46 3 Vdd
rlabel m1 33 14 33 14 3 GND
rlabel m1 33 18 33 18 3 GND
rlabel pdc 24 30 24 30 3 Vdd
rlabel m1 23 44 23 44 3 B
port 1 e
rlabel m1 23 30 23 30 3 Vdd
rlabel m1 17 33 17 33 3 Y
port 2 e
rlabel pc 20 44 20 44 3 B
port 1 e
rlabel m1 23 5 23 5 3 Y
port 2 e
rlabel m1 17 22 17 22 3 Y
port 2 e
rlabel m1 17 26 17 26 3 Y
port 2 e
rlabel m1 19 37 19 37 3 B
port 1 e
rlabel m1 19 44 19 44 3 B
port 1 e
rlabel m1 19 47 19 47 3 B
port 1 e
rlabel m1 13 44 13 44 3 A
port 3 e
rlabel pdc 17 30 17 30 3 Y
port 2 e
rlabel pc 10 44 10 44 3 A
port 3 e
rlabel m1 9 38 9 38 3 A
port 3 e
rlabel m1 9 44 9 44 3 A
port 3 e
rlabel m1 9 47 9 47 3 A
port 3 e
rlabel m1 7 30 7 30 3 Vdd
rlabel m1 7 31 7 31 3 Vdd
rlabel m1 7 34 7 34 3 Vdd
rlabel m2 30 43 30 43 3 Vdd
rlabel m2 36 15 36 15 3 GND
rlabel m2c 27 43 27 43 3 Vdd
rlabel m2c 33 15 33 15 3 GND
rlabel m2 26 35 26 35 3 Vdd
rlabel m2 26 43 26 43 3 Vdd
rlabel m2 26 46 26 46 3 Vdd
rlabel m2 13 15 13 15 3 GND
rlabel m2 13 31 13 31 3 Vdd
rlabel m2c 10 15 10 15 3 GND
rlabel m2c 10 31 10 31 3 Vdd
rlabel m2 9 14 9 14 3 GND
rlabel m2 9 15 9 15 3 GND
rlabel m2 9 18 9 18 3 GND
rlabel m2 9 30 9 30 3 Vdd
rlabel m2 9 31 9 31 3 Vdd
rlabel m2 9 34 9 34 3 Vdd
<< end >>
